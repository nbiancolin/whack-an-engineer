module part2(iResetn,iPlotBox,iBlack,iColour,iLoadX,iXY_Coord,iClock,oX,oY,oColour,oPlot,oDone);
   //specify input
   parameter X_SCREEN_PIXELS = 8'd160;
   parameter Y_SCREEN_PIXELS = 7'd120;
   input wire iResetn, iPlotBox, iBlack, iLoadX;
   input wire [2:0] iColour;
   input wire [6:0] iXY_Coord;
   input wire 	    iClock;
   output  [7:0] oX;       
   output  [6:0] oY;
   output  [2:0] oColour;     
   output  oPlot;       
   output  oDone;    

   helper u0(.iResetn(iResetn),.iPlotBox(iPlotBox),.iBlack(iBlack),
      .iColour(iColour), .iLoadX(iLoadX),.iXY_Coord(iXY_Coord),
      .clk(iClock),.oX(oX),.oY(oY), .oColour(oColour),
      .oPlot(oPlot),.oDone(oDone));
endmodule 

module helper(iResetn,iPlotBox,iBlack,iColour,iLoadX,iXY_Coord,clk,oX,oY,oColour,oPlot,oDone);
    parameter X_SCREEN_PIXELS = 8'd160;
    parameter Y_SCREEN_PIXELS = 7'd120;
    input iResetn, iPlotBox, iBlack, iLoadX;
    input [2:0] iColour;
    input [6:0] iXY_Coord;
    input clk;
    output reg [7:0] oX;      //transformed coordinates 
    output reg [6:0] oY;
    output reg [2:0] oColour;     
    output reg oPlot;       
    output reg oDone;  


    localparam  RESET        = 3'd0,
                LOADING      = 3'd1,
                DRAW_GAME    = 3'd2,
                PLOT         = 3'd3
                G_STEADY     = 3'd4,
                G_HIT        = 3'd5,
                G_RESET      = 3'd6;
    
    reg [2:0] curState, nextState;
    reg [7:0] Xsize;            //upper bound of counter
    reg [6:0] Ysize;
    reg [7:0] xProgress;        //counter
    reg [6:0] yProgress;

    reg [2:0] oColour;

    reg [15:0] counter;

    reg [1:0] selector; //used to select colours
    

    /*
    (RESET) -> reset all variables
    (LOADING) -> Clears screen (minus tape measure)
                                                                                (out) (DRAW_GAME) -> draws full game screen
    (PLOT) -> Does the plotting
    (G_STEADY) -> waits for one of 3 buttons to go to next state
    (G_HIT) -> draws the hat that has been hit
    (G_RESET) -> Draws hat back to original

    iBlack = start

    iLoadX = hit1
    iPlotBox = hit2
    iResetn = resetn


    Selector:
    00 - draw base screen
    01 - draw hh splash
    10 - draw hh outline
    */

    always@(*) begin
        case(curState)
        RESET: begin
            if(iBlack) nextState <= LOADING;
            //nextState <= iBlack ? LOADING ? RESET;
        end
        LOADING: 
            nextState <= oDone ? LOADING : PLOT;
        //DRAW_GAME:
            //nextState <= oDone ? G_STEADY : DRAW_GAME;
        //    nextState <= oDone ? LOADING: PLOT; //switches when nextState is released
        PLOT:
            nextState <= oDone ? G_STEADY : PLOT;
        G_STEADY: begin
            if(iLoadX) nextState <= G_HIT;
            else if (iPlotBox) nextState <= G_HIT;
            else if(iResetn) nextState <= RESET;
        end
        G_HIT:   
            nextState = iPlotBox ? G_HIT : PLOT; //switches on negedge
        G_RESET: 
            nextState = oDone ? G_STEADY : G_RESET;
        endcase
    end

    always@(posedge clk) begin
        if(!iResetn) curState <= RESET;
        else curState <= nextState;

        if(curState == LOADING) begin //do something
            //drawing full screen so
            oDone <= 0;
            oPlot <= 1;  
            //oColour <= 3'b000; 
            Xsize <= X_SCREEN_PIXELS - 1;
            Ysize <= Y_SCREEN_PIXELS - 1;  
            oX <= 0;
            oY <= 0;
            xProgress <= 0;
            yProgress <= 0;
            selector <= 2'b00
        end else
        //else if (curState == DRAW_GAME) begin

        //end else
        if(curState = PLOT) begin
            if (!oDone) begin
                oPlot <= 1;  
                //oColour <= oColour; 
                if (xProgress < Xsize) begin
                    oX <= oX + 1; 
                    xProgress <= xProgress + 1;  
                end else begin
                //if (xProgress == Xsize) begin
                    oX <= oX - xProgress;  
                    xProgress <= 0; 
                    if (yProgress < Ysize) begin
                        oY <= oY + 1;  
                        yProgress <= yProgress + 1; 
                    end
                end
                if (xProgress == Xsize && yProgress == Ysize) begin
                    oDone <= 1;  
                    oPlot <= 0;  
                    xSize <= 29; //xSize is for upper bound (these are now being set for hard-hat)
                    ySize <= 19;
                end
                //oColours from python script go here
                //use switch // if statements to select which colour set
                if(selector == 2'b00) begin
                    if(xProgress == 0 and yProgress == 0) oColour <= 3'b000;
                    if(xProgress == 56 and yProgress == 13) oColour <= 3'b111;
                    if(xProgress == 63 and yProgress == 13) oColour <= 3'b000;
                    if(xProgress == 55 and yProgress == 14) oColour <= 3'b111;
                    if(xProgress == 67 and yProgress == 14) oColour <= 3'b000;
                    if(xProgress == 53 and yProgress == 15) oColour <= 3'b111;
                    if(xProgress == 57 and yProgress == 15) oColour <= 3'b100;
                    if(xProgress == 62 and yProgress == 15) oColour <= 3'b111;
                    if(xProgress == 68 and yProgress == 15) oColour <= 3'b000;
                    if(xProgress == 52 and yProgress == 16) oColour <= 3'b111;
                    if(xProgress == 56 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 58 and yProgress == 16) oColour <= 3'b110;
                    if(xProgress == 61 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 66 and yProgress == 16) oColour <= 3'b111;
                    if(xProgress == 69 and yProgress == 16) oColour <= 3'b000;
                    if(xProgress == 51 and yProgress == 17) oColour <= 3'b111;
                    if(xProgress == 54 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 56 and yProgress == 17) oColour <= 3'b110;
                    if(xProgress == 57 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 58 and yProgress == 17) oColour <= 3'b110;
                    if(xProgress == 62 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 63 and yProgress == 17) oColour <= 3'b110;
                    if(xProgress == 65 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 67 and yProgress == 17) oColour <= 3'b111;
                    if(xProgress == 69 and yProgress == 17) oColour <= 3'b000;
                    if(xProgress == 50 and yProgress == 18) oColour <= 3'b111;
                    if(xProgress == 53 and yProgress == 18) oColour <= 3'b100;
                    if(xProgress == 55 and yProgress == 18) oColour <= 3'b110;
                    if(xProgress == 56 and yProgress == 18) oColour <= 3'b100;
                    if(xProgress == 57 and yProgress == 18) oColour <= 3'b110;
                    if(xProgress == 58 and yProgress == 18) oColour <= 3'b100;
                    if(xProgress == 60 and yProgress == 18) oColour <= 3'b110;
                    if(xProgress == 63 and yProgress == 18) oColour <= 3'b100;
                    if(xProgress == 65 and yProgress == 18) oColour <= 3'b110;
                    if(xProgress == 66 and yProgress == 18) oColour <= 3'b100;
                    if(xProgress == 67 and yProgress == 18) oColour <= 3'b111;
                    if(xProgress == 70 and yProgress == 18) oColour <= 3'b000;
                    if(xProgress == 49 and yProgress == 19) oColour <= 3'b111;
                    if(xProgress == 52 and yProgress == 19) oColour <= 3'b100;
                    if(xProgress == 56 and yProgress == 19) oColour <= 3'b110;
                    if(xProgress == 57 and yProgress == 19) oColour <= 3'b111;
                    if(xProgress == 58 and yProgress == 19) oColour <= 3'b110;
                    if(xProgress == 59 and yProgress == 19) oColour <= 3'b100;
                    if(xProgress == 61 and yProgress == 19) oColour <= 3'b110;
                    if(xProgress == 64 and yProgress == 19) oColour <= 3'b100;
                    if(xProgress == 68 and yProgress == 19) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 19) oColour <= 3'b000;
                    if(xProgress == 49 and yProgress == 20) oColour <= 3'b111;
                    if(xProgress == 52 and yProgress == 20) oColour <= 3'b100;
                    if(xProgress == 53 and yProgress == 20) oColour <= 3'b110;
                    if(xProgress == 55 and yProgress == 20) oColour <= 3'b111;
                    if(xProgress == 57 and yProgress == 20) oColour <= 3'b110;
                    if(xProgress == 61 and yProgress == 20) oColour <= 3'b100;
                    if(xProgress == 62 and yProgress == 20) oColour <= 3'b110;
                    if(xProgress == 65 and yProgress == 20) oColour <= 3'b100;
                    if(xProgress == 66 and yProgress == 20) oColour <= 3'b110;
                    if(xProgress == 68 and yProgress == 20) oColour <= 3'b100;
                    if(xProgress == 69 and yProgress == 20) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 20) oColour <= 3'b000;
                    if(xProgress == 49 and yProgress == 21) oColour <= 3'b111;
                    if(xProgress == 51 and yProgress == 21) oColour <= 3'b100;
                    if(xProgress == 53 and yProgress == 21) oColour <= 3'b110;
                    if(xProgress == 54 and yProgress == 21) oColour <= 3'b111;
                    if(xProgress == 56 and yProgress == 21) oColour <= 3'b110;
                    if(xProgress == 61 and yProgress == 21) oColour <= 3'b100;
                    if(xProgress == 63 and yProgress == 21) oColour <= 3'b110;
                    if(xProgress == 65 and yProgress == 21) oColour <= 3'b100;
                    if(xProgress == 67 and yProgress == 21) oColour <= 3'b110;
                    if(xProgress == 68 and yProgress == 21) oColour <= 3'b100;
                    if(xProgress == 69 and yProgress == 21) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 21) oColour <= 3'b000;
                    if(xProgress == 49 and yProgress == 22) oColour <= 3'b111;
                    if(xProgress == 51 and yProgress == 22) oColour <= 3'b100;
                    if(xProgress == 52 and yProgress == 22) oColour <= 3'b110;
                    if(xProgress == 54 and yProgress == 22) oColour <= 3'b111;
                    if(xProgress == 55 and yProgress == 22) oColour <= 3'b110;
                    if(xProgress == 62 and yProgress == 22) oColour <= 3'b100;
                    if(xProgress == 63 and yProgress == 22) oColour <= 3'b110;
                    if(xProgress == 66 and yProgress == 22) oColour <= 3'b100;
                    if(xProgress == 67 and yProgress == 22) oColour <= 3'b110;
                    if(xProgress == 69 and yProgress == 22) oColour <= 3'b100;
                    if(xProgress == 70 and yProgress == 22) oColour <= 3'b111;
                    if(xProgress == 73 and yProgress == 22) oColour <= 3'b000;
                    if(xProgress == 48 and yProgress == 23) oColour <= 3'b111;
                    if(xProgress == 51 and yProgress == 23) oColour <= 3'b100;
                    if(xProgress == 52 and yProgress == 23) oColour <= 3'b110;
                    if(xProgress == 57 and yProgress == 23) oColour <= 3'b100;
                    if(xProgress == 60 and yProgress == 23) oColour <= 3'b110;
                    if(xProgress == 62 and yProgress == 23) oColour <= 3'b100;
                    if(xProgress == 63 and yProgress == 23) oColour <= 3'b110;
                    if(xProgress == 66 and yProgress == 23) oColour <= 3'b100;
                    if(xProgress == 68 and yProgress == 23) oColour <= 3'b110;
                    if(xProgress == 69 and yProgress == 23) oColour <= 3'b100;
                    if(xProgress == 70 and yProgress == 23) oColour <= 3'b111;
                    if(xProgress == 74 and yProgress == 23) oColour <= 3'b000;
                    if(xProgress == 47 and yProgress == 24) oColour <= 3'b111;
                    if(xProgress == 50 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 52 and yProgress == 24) oColour <= 3'b110;
                    if(xProgress == 56 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 58 and yProgress == 24) oColour <= 3'b110;
                    if(xProgress == 59 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 60 and yProgress == 24) oColour <= 3'b110;
                    if(xProgress == 62 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 64 and yProgress == 24) oColour <= 3'b110;
                    if(xProgress == 67 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 68 and yProgress == 24) oColour <= 3'b110;
                    if(xProgress == 69 and yProgress == 24) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 24) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 24) oColour <= 3'b000;
                    if(xProgress == 47 and yProgress == 25) oColour <= 3'b111;
                    if(xProgress == 49 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 50 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 51 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 52 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 53 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 55 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 56 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 57 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 59 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 60 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 63 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 64 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 67 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 68 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 69 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 70 and yProgress == 25) oColour <= 3'b110;
                    if(xProgress == 71 and yProgress == 25) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 25) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 25) oColour <= 3'b000;
                    if(xProgress == 47 and yProgress == 26) oColour <= 3'b111;
                    if(xProgress == 49 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 50 and yProgress == 26) oColour <= 3'b110;
                    if(xProgress == 51 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 53 and yProgress == 26) oColour <= 3'b110;
                    if(xProgress == 55 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 60 and yProgress == 26) oColour <= 3'b110;
                    if(xProgress == 63 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 64 and yProgress == 26) oColour <= 3'b110;
                    if(xProgress == 67 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 69 and yProgress == 26) oColour <= 3'b110;
                    if(xProgress == 72 and yProgress == 26) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 26) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 26) oColour <= 3'b000;
                    if(xProgress == 47 and yProgress == 27) oColour <= 3'b111;
                    if(xProgress == 50 and yProgress == 27) oColour <= 3'b100;
                    if(xProgress == 51 and yProgress == 27) oColour <= 3'b110;
                    if(xProgress == 53 and yProgress == 27) oColour <= 3'b100;
                    if(xProgress == 55 and yProgress == 27) oColour <= 3'b110;
                    if(xProgress == 57 and yProgress == 27) oColour <= 3'b100;
                    if(xProgress == 59 and yProgress == 27) oColour <= 3'b110;
                    if(xProgress == 60 and yProgress == 27) oColour <= 3'b100;
                    if(xProgress == 68 and yProgress == 27) oColour <= 3'b110;
                    if(xProgress == 72 and yProgress == 27) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 27) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 27) oColour <= 3'b000;
                    if(xProgress == 48 and yProgress == 28) oColour <= 3'b111;
                    if(xProgress == 51 and yProgress == 28) oColour <= 3'b100;
                    if(xProgress == 55 and yProgress == 28) oColour <= 3'b110;
                    if(xProgress == 71 and yProgress == 28) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 28) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 28) oColour <= 3'b000;
                    if(xProgress == 49 and yProgress == 29) oColour <= 3'b111;
                    if(xProgress == 54 and yProgress == 29) oColour <= 3'b100;
                    if(xProgress == 57 and yProgress == 29) oColour <= 3'b110;
                    if(xProgress == 70 and yProgress == 29) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 29) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 29) oColour <= 3'b000;
                    if(xProgress == 50 and yProgress == 30) oColour <= 3'b111;
                    if(xProgress == 56 and yProgress == 30) oColour <= 3'b100;
                    if(xProgress == 71 and yProgress == 30) oColour <= 3'b111;
                    if(xProgress == 74 and yProgress == 30) oColour <= 3'b000;
                    if(xProgress == 53 and yProgress == 31) oColour <= 3'b111;
                    if(xProgress == 73 and yProgress == 31) oColour <= 3'b000;
                    if(xProgress == 106 and yProgress == 31) oColour <= 3'b111;
                    if(xProgress == 113 and yProgress == 31) oColour <= 3'b000;
                    if(xProgress == 55 and yProgress == 32) oColour <= 3'b111;
                    if(xProgress == 72 and yProgress == 32) oColour <= 3'b000;
                    if(xProgress == 105 and yProgress == 32) oColour <= 3'b111;
                    if(xProgress == 117 and yProgress == 32) oColour <= 3'b000;
                    if(xProgress == 103 and yProgress == 33) oColour <= 3'b111;
                    if(xProgress == 107 and yProgress == 33) oColour <= 3'b100;
                    if(xProgress == 112 and yProgress == 33) oColour <= 3'b111;
                    if(xProgress == 118 and yProgress == 33) oColour <= 3'b000;
                    if(xProgress == 102 and yProgress == 34) oColour <= 3'b111;
                    if(xProgress == 106 and yProgress == 34) oColour <= 3'b100;
                    if(xProgress == 108 and yProgress == 34) oColour <= 3'b110;
                    if(xProgress == 111 and yProgress == 34) oColour <= 3'b100;
                    if(xProgress == 116 and yProgress == 34) oColour <= 3'b111;
                    if(xProgress == 119 and yProgress == 34) oColour <= 3'b000;
                    if(xProgress == 101 and yProgress == 35) oColour <= 3'b111;
                    if(xProgress == 104 and yProgress == 35) oColour <= 3'b100;
                    if(xProgress == 106 and yProgress == 35) oColour <= 3'b110;
                    if(xProgress == 107 and yProgress == 35) oColour <= 3'b100;
                    if(xProgress == 108 and yProgress == 35) oColour <= 3'b110;
                    if(xProgress == 112 and yProgress == 35) oColour <= 3'b100;
                    if(xProgress == 113 and yProgress == 35) oColour <= 3'b110;
                    if(xProgress == 115 and yProgress == 35) oColour <= 3'b100;
                    if(xProgress == 117 and yProgress == 35) oColour <= 3'b111;
                    if(xProgress == 119 and yProgress == 35) oColour <= 3'b000;
                    if(xProgress == 100 and yProgress == 36) oColour <= 3'b111;
                    if(xProgress == 103 and yProgress == 36) oColour <= 3'b100;
                    if(xProgress == 105 and yProgress == 36) oColour <= 3'b110;
                    if(xProgress == 106 and yProgress == 36) oColour <= 3'b100;
                    if(xProgress == 107 and yProgress == 36) oColour <= 3'b110;
                    if(xProgress == 108 and yProgress == 36) oColour <= 3'b100;
                    if(xProgress == 110 and yProgress == 36) oColour <= 3'b110;
                    if(xProgress == 113 and yProgress == 36) oColour <= 3'b100;
                    if(xProgress == 115 and yProgress == 36) oColour <= 3'b110;
                    if(xProgress == 116 and yProgress == 36) oColour <= 3'b100;
                    if(xProgress == 117 and yProgress == 36) oColour <= 3'b111;
                    if(xProgress == 120 and yProgress == 36) oColour <= 3'b000;
                    if(xProgress == 99 and yProgress == 37) oColour <= 3'b111;
                    if(xProgress == 102 and yProgress == 37) oColour <= 3'b100;
                    if(xProgress == 106 and yProgress == 37) oColour <= 3'b110;
                    if(xProgress == 107 and yProgress == 37) oColour <= 3'b111;
                    if(xProgress == 108 and yProgress == 37) oColour <= 3'b110;
                    if(xProgress == 109 and yProgress == 37) oColour <= 3'b100;
                    if(xProgress == 111 and yProgress == 37) oColour <= 3'b110;
                    if(xProgress == 114 and yProgress == 37) oColour <= 3'b100;
                    if(xProgress == 118 and yProgress == 37) oColour <= 3'b111;
                    if(xProgress == 121 and yProgress == 37) oColour <= 3'b000;
                    if(xProgress == 99 and yProgress == 38) oColour <= 3'b111;
                    if(xProgress == 102 and yProgress == 38) oColour <= 3'b100;
                    if(xProgress == 103 and yProgress == 38) oColour <= 3'b110;
                    if(xProgress == 105 and yProgress == 38) oColour <= 3'b111;
                    if(xProgress == 107 and yProgress == 38) oColour <= 3'b110;
                    if(xProgress == 111 and yProgress == 38) oColour <= 3'b100;
                    if(xProgress == 112 and yProgress == 38) oColour <= 3'b110;
                    if(xProgress == 115 and yProgress == 38) oColour <= 3'b100;
                    if(xProgress == 116 and yProgress == 38) oColour <= 3'b110;
                    if(xProgress == 118 and yProgress == 38) oColour <= 3'b100;
                    if(xProgress == 119 and yProgress == 38) oColour <= 3'b111;
                    if(xProgress == 121 and yProgress == 38) oColour <= 3'b000;
                    if(xProgress == 99 and yProgress == 39) oColour <= 3'b111;
                    if(xProgress == 101 and yProgress == 39) oColour <= 3'b100;
                    if(xProgress == 103 and yProgress == 39) oColour <= 3'b110;
                    if(xProgress == 104 and yProgress == 39) oColour <= 3'b111;
                    if(xProgress == 106 and yProgress == 39) oColour <= 3'b110;
                    if(xProgress == 111 and yProgress == 39) oColour <= 3'b100;
                    if(xProgress == 113 and yProgress == 39) oColour <= 3'b110;
                    if(xProgress == 115 and yProgress == 39) oColour <= 3'b100;
                    if(xProgress == 117 and yProgress == 39) oColour <= 3'b110;
                    if(xProgress == 118 and yProgress == 39) oColour <= 3'b100;
                    if(xProgress == 119 and yProgress == 39) oColour <= 3'b111;
                    if(xProgress == 121 and yProgress == 39) oColour <= 3'b000;
                    if(xProgress == 99 and yProgress == 40) oColour <= 3'b111;
                    if(xProgress == 101 and yProgress == 40) oColour <= 3'b100;
                    if(xProgress == 102 and yProgress == 40) oColour <= 3'b110;
                    if(xProgress == 104 and yProgress == 40) oColour <= 3'b111;
                    if(xProgress == 105 and yProgress == 40) oColour <= 3'b110;
                    if(xProgress == 112 and yProgress == 40) oColour <= 3'b100;
                    if(xProgress == 113 and yProgress == 40) oColour <= 3'b110;
                    if(xProgress == 116 and yProgress == 40) oColour <= 3'b100;
                    if(xProgress == 117 and yProgress == 40) oColour <= 3'b110;
                    if(xProgress == 119 and yProgress == 40) oColour <= 3'b100;
                    if(xProgress == 120 and yProgress == 40) oColour <= 3'b111;
                    if(xProgress == 123 and yProgress == 40) oColour <= 3'b000;
                    if(xProgress == 98 and yProgress == 41) oColour <= 3'b111;
                    if(xProgress == 101 and yProgress == 41) oColour <= 3'b100;
                    if(xProgress == 102 and yProgress == 41) oColour <= 3'b110;
                    if(xProgress == 107 and yProgress == 41) oColour <= 3'b100;
                    if(xProgress == 110 and yProgress == 41) oColour <= 3'b110;
                    if(xProgress == 112 and yProgress == 41) oColour <= 3'b100;
                    if(xProgress == 113 and yProgress == 41) oColour <= 3'b110;
                    if(xProgress == 116 and yProgress == 41) oColour <= 3'b100;
                    if(xProgress == 118 and yProgress == 41) oColour <= 3'b110;
                    if(xProgress == 119 and yProgress == 41) oColour <= 3'b100;
                    if(xProgress == 120 and yProgress == 41) oColour <= 3'b111;
                    if(xProgress == 124 and yProgress == 41) oColour <= 3'b000;
                    if(xProgress == 97 and yProgress == 42) oColour <= 3'b111;
                    if(xProgress == 100 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 102 and yProgress == 42) oColour <= 3'b110;
                    if(xProgress == 106 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 108 and yProgress == 42) oColour <= 3'b110;
                    if(xProgress == 109 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 110 and yProgress == 42) oColour <= 3'b110;
                    if(xProgress == 112 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 114 and yProgress == 42) oColour <= 3'b110;
                    if(xProgress == 117 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 118 and yProgress == 42) oColour <= 3'b110;
                    if(xProgress == 119 and yProgress == 42) oColour <= 3'b100;
                    if(xProgress == 122 and yProgress == 42) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 42) oColour <= 3'b000;
                    if(xProgress == 97 and yProgress == 43) oColour <= 3'b111;
                    if(xProgress == 99 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 100 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 101 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 102 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 103 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 105 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 106 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 107 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 109 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 110 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 113 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 114 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 117 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 118 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 119 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 120 and yProgress == 43) oColour <= 3'b110;
                    if(xProgress == 121 and yProgress == 43) oColour <= 3'b100;
                    if(xProgress == 123 and yProgress == 43) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 43) oColour <= 3'b000;
                    if(xProgress == 97 and yProgress == 44) oColour <= 3'b111;
                    if(xProgress == 99 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 100 and yProgress == 44) oColour <= 3'b110;
                    if(xProgress == 101 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 103 and yProgress == 44) oColour <= 3'b110;
                    if(xProgress == 105 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 110 and yProgress == 44) oColour <= 3'b110;
                    if(xProgress == 113 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 114 and yProgress == 44) oColour <= 3'b110;
                    if(xProgress == 117 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 119 and yProgress == 44) oColour <= 3'b110;
                    if(xProgress == 122 and yProgress == 44) oColour <= 3'b100;
                    if(xProgress == 123 and yProgress == 44) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 44) oColour <= 3'b000;
                    if(xProgress == 97 and yProgress == 45) oColour <= 3'b111;
                    if(xProgress == 100 and yProgress == 45) oColour <= 3'b100;
                    if(xProgress == 101 and yProgress == 45) oColour <= 3'b110;
                    if(xProgress == 103 and yProgress == 45) oColour <= 3'b100;
                    if(xProgress == 105 and yProgress == 45) oColour <= 3'b110;
                    if(xProgress == 107 and yProgress == 45) oColour <= 3'b100;
                    if(xProgress == 109 and yProgress == 45) oColour <= 3'b110;
                    if(xProgress == 110 and yProgress == 45) oColour <= 3'b100;
                    if(xProgress == 118 and yProgress == 45) oColour <= 3'b110;
                    if(xProgress == 122 and yProgress == 45) oColour <= 3'b100;
                    if(xProgress == 123 and yProgress == 45) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 45) oColour <= 3'b000;
                    if(xProgress == 98 and yProgress == 46) oColour <= 3'b111;
                    if(xProgress == 101 and yProgress == 46) oColour <= 3'b100;
                    if(xProgress == 105 and yProgress == 46) oColour <= 3'b110;
                    if(xProgress == 121 and yProgress == 46) oColour <= 3'b100;
                    if(xProgress == 123 and yProgress == 46) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 46) oColour <= 3'b000;
                    if(xProgress == 99 and yProgress == 47) oColour <= 3'b111;
                    if(xProgress == 104 and yProgress == 47) oColour <= 3'b100;
                    if(xProgress == 107 and yProgress == 47) oColour <= 3'b110;
                    if(xProgress == 120 and yProgress == 47) oColour <= 3'b100;
                    if(xProgress == 122 and yProgress == 47) oColour <= 3'b111;
                    if(xProgress == 125 and yProgress == 47) oColour <= 3'b000;
                    if(xProgress == 100 and yProgress == 48) oColour <= 3'b111;
                    if(xProgress == 106 and yProgress == 48) oColour <= 3'b100;
                    if(xProgress == 121 and yProgress == 48) oColour <= 3'b111;
                    if(xProgress == 124 and yProgress == 48) oColour <= 3'b000;
                    if(xProgress == 103 and yProgress == 49) oColour <= 3'b111;
                    if(xProgress == 123 and yProgress == 49) oColour <= 3'b000;
                    if(xProgress == 105 and yProgress == 50) oColour <= 3'b111;
                    if(xProgress == 122 and yProgress == 50) oColour <= 3'b000;
                    if(xProgress == 19 and yProgress == 53) oColour <= 3'b111;
                    if(xProgress == 26 and yProgress == 53) oColour <= 3'b000;
                    if(xProgress == 18 and yProgress == 54) oColour <= 3'b111;
                    if(xProgress == 30 and yProgress == 54) oColour <= 3'b000;
                    if(xProgress == 16 and yProgress == 55) oColour <= 3'b111;
                    if(xProgress == 20 and yProgress == 55) oColour <= 3'b100;
                    if(xProgress == 25 and yProgress == 55) oColour <= 3'b111;
                    if(xProgress == 31 and yProgress == 55) oColour <= 3'b000;
                    if(xProgress == 15 and yProgress == 56) oColour <= 3'b111;
                    if(xProgress == 19 and yProgress == 56) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 56) oColour <= 3'b110;
                    if(xProgress == 24 and yProgress == 56) oColour <= 3'b100;
                    if(xProgress == 29 and yProgress == 56) oColour <= 3'b111;
                    if(xProgress == 32 and yProgress == 56) oColour <= 3'b000;
                    if(xProgress == 14 and yProgress == 57) oColour <= 3'b111;
                    if(xProgress == 17 and yProgress == 57) oColour <= 3'b100;
                    if(xProgress == 19 and yProgress == 57) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 57) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 57) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 57) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 57) oColour <= 3'b110;
                    if(xProgress == 28 and yProgress == 57) oColour <= 3'b100;
                    if(xProgress == 30 and yProgress == 57) oColour <= 3'b111;
                    if(xProgress == 32 and yProgress == 57) oColour <= 3'b000;
                    if(xProgress == 13 and yProgress == 58) oColour <= 3'b111;
                    if(xProgress == 16 and yProgress == 58) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 58) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 58) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 58) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 58) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 58) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 58) oColour <= 3'b100;
                    if(xProgress == 28 and yProgress == 58) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 58) oColour <= 3'b100;
                    if(xProgress == 30 and yProgress == 58) oColour <= 3'b111;
                    if(xProgress == 33 and yProgress == 58) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 59) oColour <= 3'b111;
                    if(xProgress == 15 and yProgress == 59) oColour <= 3'b100;
                    if(xProgress == 19 and yProgress == 59) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 59) oColour <= 3'b111;
                    if(xProgress == 21 and yProgress == 59) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 59) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 59) oColour <= 3'b110;
                    if(xProgress == 27 and yProgress == 59) oColour <= 3'b100;
                    if(xProgress == 31 and yProgress == 59) oColour <= 3'b111;
                    if(xProgress == 34 and yProgress == 59) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 60) oColour <= 3'b111;
                    if(xProgress == 15 and yProgress == 60) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 60) oColour <= 3'b110;
                    if(xProgress == 18 and yProgress == 60) oColour <= 3'b111;
                    if(xProgress == 20 and yProgress == 60) oColour <= 3'b110;
                    if(xProgress == 24 and yProgress == 60) oColour <= 3'b100;
                    if(xProgress == 25 and yProgress == 60) oColour <= 3'b110;
                    if(xProgress == 28 and yProgress == 60) oColour <= 3'b100;
                    if(xProgress == 29 and yProgress == 60) oColour <= 3'b110;
                    if(xProgress == 31 and yProgress == 60) oColour <= 3'b100;
                    if(xProgress == 32 and yProgress == 60) oColour <= 3'b111;
                    if(xProgress == 34 and yProgress == 60) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 61) oColour <= 3'b111;
                    if(xProgress == 14 and yProgress == 61) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 61) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 61) oColour <= 3'b111;
                    if(xProgress == 19 and yProgress == 61) oColour <= 3'b110;
                    if(xProgress == 24 and yProgress == 61) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 61) oColour <= 3'b110;
                    if(xProgress == 28 and yProgress == 61) oColour <= 3'b100;
                    if(xProgress == 30 and yProgress == 61) oColour <= 3'b110;
                    if(xProgress == 31 and yProgress == 61) oColour <= 3'b100;
                    if(xProgress == 32 and yProgress == 61) oColour <= 3'b111;
                    if(xProgress == 34 and yProgress == 61) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 62) oColour <= 3'b111;
                    if(xProgress == 14 and yProgress == 62) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 62) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 62) oColour <= 3'b111;
                    if(xProgress == 18 and yProgress == 62) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 62) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 62) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 62) oColour <= 3'b100;
                    if(xProgress == 30 and yProgress == 62) oColour <= 3'b110;
                    if(xProgress == 32 and yProgress == 62) oColour <= 3'b100;
                    if(xProgress == 33 and yProgress == 62) oColour <= 3'b111;
                    if(xProgress == 36 and yProgress == 62) oColour <= 3'b000;
                    if(xProgress == 11 and yProgress == 63) oColour <= 3'b111;
                    if(xProgress == 14 and yProgress == 63) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 63) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 63) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 63) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 63) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 63) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 63) oColour <= 3'b100;
                    if(xProgress == 31 and yProgress == 63) oColour <= 3'b110;
                    if(xProgress == 32 and yProgress == 63) oColour <= 3'b100;
                    if(xProgress == 33 and yProgress == 63) oColour <= 3'b111;
                    if(xProgress == 37 and yProgress == 63) oColour <= 3'b000;
                    if(xProgress == 135 and yProgress == 63) oColour <= 3'b111;
                    if(xProgress == 142 and yProgress == 63) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 64) oColour <= 3'b111;
                    if(xProgress == 13 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 64) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 64) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 64) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 64) oColour <= 3'b110;
                    if(xProgress == 30 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 31 and yProgress == 64) oColour <= 3'b110;
                    if(xProgress == 32 and yProgress == 64) oColour <= 3'b100;
                    if(xProgress == 35 and yProgress == 64) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 64) oColour <= 3'b000;
                    if(xProgress == 134 and yProgress == 64) oColour <= 3'b111;
                    if(xProgress == 146 and yProgress == 64) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 65) oColour <= 3'b111;
                    if(xProgress == 12 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 13 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 14 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 30 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 31 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 32 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 33 and yProgress == 65) oColour <= 3'b110;
                    if(xProgress == 34 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 36 and yProgress == 65) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 65) oColour <= 3'b000;
                    if(xProgress == 132 and yProgress == 65) oColour <= 3'b111;
                    if(xProgress == 136 and yProgress == 65) oColour <= 3'b100;
                    if(xProgress == 141 and yProgress == 65) oColour <= 3'b111;
                    if(xProgress == 147 and yProgress == 65) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 66) oColour <= 3'b111;
                    if(xProgress == 12 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 13 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 14 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 18 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 30 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 32 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 35 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 36 and yProgress == 66) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 66) oColour <= 3'b000;
                    if(xProgress == 131 and yProgress == 66) oColour <= 3'b111;
                    if(xProgress == 135 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 137 and yProgress == 66) oColour <= 3'b110;
                    if(xProgress == 140 and yProgress == 66) oColour <= 3'b100;
                    if(xProgress == 145 and yProgress == 66) oColour <= 3'b111;
                    if(xProgress == 148 and yProgress == 66) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 67) oColour <= 3'b111;
                    if(xProgress == 13 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 31 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 35 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 36 and yProgress == 67) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 67) oColour <= 3'b000;
                    if(xProgress == 130 and yProgress == 67) oColour <= 3'b111;
                    if(xProgress == 133 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 135 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 136 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 137 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 141 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 142 and yProgress == 67) oColour <= 3'b110;
                    if(xProgress == 144 and yProgress == 67) oColour <= 3'b100;
                    if(xProgress == 146 and yProgress == 67) oColour <= 3'b111;
                    if(xProgress == 148 and yProgress == 67) oColour <= 3'b000;
                    if(xProgress == 11 and yProgress == 68) oColour <= 3'b111;
                    if(xProgress == 14 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 68) oColour <= 3'b110;
                    if(xProgress == 34 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 36 and yProgress == 68) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 68) oColour <= 3'b000;
                    if(xProgress == 129 and yProgress == 68) oColour <= 3'b111;
                    if(xProgress == 132 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 134 and yProgress == 68) oColour <= 3'b110;
                    if(xProgress == 135 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 136 and yProgress == 68) oColour <= 3'b110;
                    if(xProgress == 137 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 139 and yProgress == 68) oColour <= 3'b110;
                    if(xProgress == 142 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 144 and yProgress == 68) oColour <= 3'b110;
                    if(xProgress == 145 and yProgress == 68) oColour <= 3'b100;
                    if(xProgress == 146 and yProgress == 68) oColour <= 3'b111;
                    if(xProgress == 149 and yProgress == 68) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 69) oColour <= 3'b111;
                    if(xProgress == 17 and yProgress == 69) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 69) oColour <= 3'b110;
                    if(xProgress == 33 and yProgress == 69) oColour <= 3'b100;
                    if(xProgress == 35 and yProgress == 69) oColour <= 3'b111;
                    if(xProgress == 38 and yProgress == 69) oColour <= 3'b000;
                    if(xProgress == 128 and yProgress == 69) oColour <= 3'b111;
                    if(xProgress == 131 and yProgress == 69) oColour <= 3'b100;
                    if(xProgress == 135 and yProgress == 69) oColour <= 3'b110;
                    if(xProgress == 136 and yProgress == 69) oColour <= 3'b111;
                    if(xProgress == 137 and yProgress == 69) oColour <= 3'b110;
                    if(xProgress == 138 and yProgress == 69) oColour <= 3'b100;
                    if(xProgress == 140 and yProgress == 69) oColour <= 3'b110;
                    if(xProgress == 143 and yProgress == 69) oColour <= 3'b100;
                    if(xProgress == 147 and yProgress == 69) oColour <= 3'b111;
                    if(xProgress == 150 and yProgress == 69) oColour <= 3'b000;
                    if(xProgress == 13 and yProgress == 70) oColour <= 3'b111;
                    if(xProgress == 19 and yProgress == 70) oColour <= 3'b100;
                    if(xProgress == 34 and yProgress == 70) oColour <= 3'b111;
                    if(xProgress == 37 and yProgress == 70) oColour <= 3'b000;
                    if(xProgress == 128 and yProgress == 70) oColour <= 3'b111;
                    if(xProgress == 131 and yProgress == 70) oColour <= 3'b100;
                    if(xProgress == 132 and yProgress == 70) oColour <= 3'b110;
                    if(xProgress == 134 and yProgress == 70) oColour <= 3'b111;
                    if(xProgress == 136 and yProgress == 70) oColour <= 3'b110;
                    if(xProgress == 140 and yProgress == 70) oColour <= 3'b100;
                    if(xProgress == 141 and yProgress == 70) oColour <= 3'b110;
                    if(xProgress == 144 and yProgress == 70) oColour <= 3'b100;
                    if(xProgress == 145 and yProgress == 70) oColour <= 3'b110;
                    if(xProgress == 147 and yProgress == 70) oColour <= 3'b100;
                    if(xProgress == 148 and yProgress == 70) oColour <= 3'b111;
                    if(xProgress == 150 and yProgress == 70) oColour <= 3'b000;
                    if(xProgress == 16 and yProgress == 71) oColour <= 3'b111;
                    if(xProgress == 36 and yProgress == 71) oColour <= 3'b000;
                    if(xProgress == 128 and yProgress == 71) oColour <= 3'b111;
                    if(xProgress == 130 and yProgress == 71) oColour <= 3'b100;
                    if(xProgress == 132 and yProgress == 71) oColour <= 3'b110;
                    if(xProgress == 133 and yProgress == 71) oColour <= 3'b111;
                    if(xProgress == 135 and yProgress == 71) oColour <= 3'b110;
                    if(xProgress == 140 and yProgress == 71) oColour <= 3'b100;
                    if(xProgress == 142 and yProgress == 71) oColour <= 3'b110;
                    if(xProgress == 144 and yProgress == 71) oColour <= 3'b100;
                    if(xProgress == 146 and yProgress == 71) oColour <= 3'b110;
                    if(xProgress == 147 and yProgress == 71) oColour <= 3'b100;
                    if(xProgress == 148 and yProgress == 71) oColour <= 3'b111;
                    if(xProgress == 150 and yProgress == 71) oColour <= 3'b000;
                    if(xProgress == 18 and yProgress == 72) oColour <= 3'b111;
                    if(xProgress == 35 and yProgress == 72) oColour <= 3'b000;
                    if(xProgress == 128 and yProgress == 72) oColour <= 3'b111;
                    if(xProgress == 130 and yProgress == 72) oColour <= 3'b100;
                    if(xProgress == 131 and yProgress == 72) oColour <= 3'b110;
                    if(xProgress == 133 and yProgress == 72) oColour <= 3'b111;
                    if(xProgress == 134 and yProgress == 72) oColour <= 3'b110;
                    if(xProgress == 141 and yProgress == 72) oColour <= 3'b100;
                    if(xProgress == 142 and yProgress == 72) oColour <= 3'b110;
                    if(xProgress == 145 and yProgress == 72) oColour <= 3'b100;
                    if(xProgress == 146 and yProgress == 72) oColour <= 3'b110;
                    if(xProgress == 148 and yProgress == 72) oColour <= 3'b100;
                    if(xProgress == 149 and yProgress == 72) oColour <= 3'b111;
                    if(xProgress == 152 and yProgress == 72) oColour <= 3'b000;
                    if(xProgress == 127 and yProgress == 73) oColour <= 3'b111;
                    if(xProgress == 130 and yProgress == 73) oColour <= 3'b100;
                    if(xProgress == 131 and yProgress == 73) oColour <= 3'b110;
                    if(xProgress == 136 and yProgress == 73) oColour <= 3'b100;
                    if(xProgress == 139 and yProgress == 73) oColour <= 3'b110;
                    if(xProgress == 141 and yProgress == 73) oColour <= 3'b100;
                    if(xProgress == 142 and yProgress == 73) oColour <= 3'b110;
                    if(xProgress == 145 and yProgress == 73) oColour <= 3'b100;
                    if(xProgress == 147 and yProgress == 73) oColour <= 3'b110;
                    if(xProgress == 148 and yProgress == 73) oColour <= 3'b100;
                    if(xProgress == 149 and yProgress == 73) oColour <= 3'b111;
                    if(xProgress == 153 and yProgress == 73) oColour <= 3'b000;
                    if(xProgress == 126 and yProgress == 74) oColour <= 3'b111;
                    if(xProgress == 129 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 131 and yProgress == 74) oColour <= 3'b110;
                    if(xProgress == 135 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 137 and yProgress == 74) oColour <= 3'b110;
                    if(xProgress == 138 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 139 and yProgress == 74) oColour <= 3'b110;
                    if(xProgress == 141 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 143 and yProgress == 74) oColour <= 3'b110;
                    if(xProgress == 146 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 147 and yProgress == 74) oColour <= 3'b110;
                    if(xProgress == 148 and yProgress == 74) oColour <= 3'b100;
                    if(xProgress == 151 and yProgress == 74) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 74) oColour <= 3'b000;
                    if(xProgress == 126 and yProgress == 75) oColour <= 3'b111;
                    if(xProgress == 128 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 129 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 130 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 131 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 132 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 134 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 135 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 136 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 138 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 139 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 142 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 143 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 146 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 147 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 148 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 149 and yProgress == 75) oColour <= 3'b110;
                    if(xProgress == 150 and yProgress == 75) oColour <= 3'b100;
                    if(xProgress == 152 and yProgress == 75) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 75) oColour <= 3'b000;
                    if(xProgress == 126 and yProgress == 76) oColour <= 3'b111;
                    if(xProgress == 128 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 129 and yProgress == 76) oColour <= 3'b110;
                    if(xProgress == 130 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 132 and yProgress == 76) oColour <= 3'b110;
                    if(xProgress == 134 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 139 and yProgress == 76) oColour <= 3'b110;
                    if(xProgress == 142 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 143 and yProgress == 76) oColour <= 3'b110;
                    if(xProgress == 146 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 148 and yProgress == 76) oColour <= 3'b110;
                    if(xProgress == 151 and yProgress == 76) oColour <= 3'b100;
                    if(xProgress == 152 and yProgress == 76) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 76) oColour <= 3'b000;
                    if(xProgress == 126 and yProgress == 77) oColour <= 3'b111;
                    if(xProgress == 129 and yProgress == 77) oColour <= 3'b100;
                    if(xProgress == 130 and yProgress == 77) oColour <= 3'b110;
                    if(xProgress == 132 and yProgress == 77) oColour <= 3'b100;
                    if(xProgress == 134 and yProgress == 77) oColour <= 3'b110;
                    if(xProgress == 136 and yProgress == 77) oColour <= 3'b100;
                    if(xProgress == 138 and yProgress == 77) oColour <= 3'b110;
                    if(xProgress == 139 and yProgress == 77) oColour <= 3'b100;
                    if(xProgress == 147 and yProgress == 77) oColour <= 3'b110;
                    if(xProgress == 151 and yProgress == 77) oColour <= 3'b100;
                    if(xProgress == 152 and yProgress == 77) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 77) oColour <= 3'b000;
                    if(xProgress == 127 and yProgress == 78) oColour <= 3'b111;
                    if(xProgress == 130 and yProgress == 78) oColour <= 3'b100;
                    if(xProgress == 134 and yProgress == 78) oColour <= 3'b110;
                    if(xProgress == 150 and yProgress == 78) oColour <= 3'b100;
                    if(xProgress == 152 and yProgress == 78) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 78) oColour <= 3'b000;
                    if(xProgress == 128 and yProgress == 79) oColour <= 3'b111;
                    if(xProgress == 133 and yProgress == 79) oColour <= 3'b100;
                    if(xProgress == 136 and yProgress == 79) oColour <= 3'b110;
                    if(xProgress == 149 and yProgress == 79) oColour <= 3'b100;
                    if(xProgress == 151 and yProgress == 79) oColour <= 3'b111;
                    if(xProgress == 154 and yProgress == 79) oColour <= 3'b000;
                    if(xProgress == 129 and yProgress == 80) oColour <= 3'b111;
                    if(xProgress == 135 and yProgress == 80) oColour <= 3'b100;
                    if(xProgress == 150 and yProgress == 80) oColour <= 3'b111;
                    if(xProgress == 153 and yProgress == 80) oColour <= 3'b000;
                    if(xProgress == 132 and yProgress == 81) oColour <= 3'b111;
                    if(xProgress == 152 and yProgress == 81) oColour <= 3'b000;
                    if(xProgress == 76 and yProgress == 82) oColour <= 3'b111;
                    if(xProgress == 83 and yProgress == 82) oColour <= 3'b000;
                    if(xProgress == 134 and yProgress == 82) oColour <= 3'b111;
                    if(xProgress == 151 and yProgress == 82) oColour <= 3'b000;
                    if(xProgress == 75 and yProgress == 83) oColour <= 3'b111;
                    if(xProgress == 87 and yProgress == 83) oColour <= 3'b000;
                    if(xProgress == 73 and yProgress == 84) oColour <= 3'b111;
                    if(xProgress == 77 and yProgress == 84) oColour <= 3'b100;
                    if(xProgress == 82 and yProgress == 84) oColour <= 3'b111;
                    if(xProgress == 88 and yProgress == 84) oColour <= 3'b000;
                    if(xProgress == 72 and yProgress == 85) oColour <= 3'b111;
                    if(xProgress == 76 and yProgress == 85) oColour <= 3'b100;
                    if(xProgress == 78 and yProgress == 85) oColour <= 3'b110;
                    if(xProgress == 81 and yProgress == 85) oColour <= 3'b100;
                    if(xProgress == 86 and yProgress == 85) oColour <= 3'b111;
                    if(xProgress == 89 and yProgress == 85) oColour <= 3'b000;
                    if(xProgress == 71 and yProgress == 86) oColour <= 3'b111;
                    if(xProgress == 74 and yProgress == 86) oColour <= 3'b100;
                    if(xProgress == 76 and yProgress == 86) oColour <= 3'b110;
                    if(xProgress == 77 and yProgress == 86) oColour <= 3'b100;
                    if(xProgress == 78 and yProgress == 86) oColour <= 3'b110;
                    if(xProgress == 82 and yProgress == 86) oColour <= 3'b100;
                    if(xProgress == 83 and yProgress == 86) oColour <= 3'b110;
                    if(xProgress == 85 and yProgress == 86) oColour <= 3'b100;
                    if(xProgress == 87 and yProgress == 86) oColour <= 3'b111;
                    if(xProgress == 89 and yProgress == 86) oColour <= 3'b000;
                    if(xProgress == 70 and yProgress == 87) oColour <= 3'b111;
                    if(xProgress == 73 and yProgress == 87) oColour <= 3'b100;
                    if(xProgress == 75 and yProgress == 87) oColour <= 3'b110;
                    if(xProgress == 76 and yProgress == 87) oColour <= 3'b100;
                    if(xProgress == 77 and yProgress == 87) oColour <= 3'b110;
                    if(xProgress == 78 and yProgress == 87) oColour <= 3'b100;
                    if(xProgress == 80 and yProgress == 87) oColour <= 3'b110;
                    if(xProgress == 83 and yProgress == 87) oColour <= 3'b100;
                    if(xProgress == 85 and yProgress == 87) oColour <= 3'b110;
                    if(xProgress == 86 and yProgress == 87) oColour <= 3'b100;
                    if(xProgress == 87 and yProgress == 87) oColour <= 3'b111;
                    if(xProgress == 90 and yProgress == 87) oColour <= 3'b000;
                    if(xProgress == 69 and yProgress == 88) oColour <= 3'b111;
                    if(xProgress == 72 and yProgress == 88) oColour <= 3'b100;
                    if(xProgress == 76 and yProgress == 88) oColour <= 3'b110;
                    if(xProgress == 77 and yProgress == 88) oColour <= 3'b111;
                    if(xProgress == 78 and yProgress == 88) oColour <= 3'b110;
                    if(xProgress == 79 and yProgress == 88) oColour <= 3'b100;
                    if(xProgress == 81 and yProgress == 88) oColour <= 3'b110;
                    if(xProgress == 84 and yProgress == 88) oColour <= 3'b100;
                    if(xProgress == 88 and yProgress == 88) oColour <= 3'b111;
                    if(xProgress == 91 and yProgress == 88) oColour <= 3'b000;
                    if(xProgress == 69 and yProgress == 89) oColour <= 3'b111;
                    if(xProgress == 72 and yProgress == 89) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 89) oColour <= 3'b110;
                    if(xProgress == 75 and yProgress == 89) oColour <= 3'b111;
                    if(xProgress == 77 and yProgress == 89) oColour <= 3'b110;
                    if(xProgress == 81 and yProgress == 89) oColour <= 3'b100;
                    if(xProgress == 82 and yProgress == 89) oColour <= 3'b110;
                    if(xProgress == 85 and yProgress == 89) oColour <= 3'b100;
                    if(xProgress == 86 and yProgress == 89) oColour <= 3'b110;
                    if(xProgress == 88 and yProgress == 89) oColour <= 3'b100;
                    if(xProgress == 89 and yProgress == 89) oColour <= 3'b111;
                    if(xProgress == 91 and yProgress == 89) oColour <= 3'b000;
                    if(xProgress == 69 and yProgress == 90) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 90) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 90) oColour <= 3'b110;
                    if(xProgress == 74 and yProgress == 90) oColour <= 3'b111;
                    if(xProgress == 76 and yProgress == 90) oColour <= 3'b110;
                    if(xProgress == 81 and yProgress == 90) oColour <= 3'b100;
                    if(xProgress == 83 and yProgress == 90) oColour <= 3'b110;
                    if(xProgress == 85 and yProgress == 90) oColour <= 3'b100;
                    if(xProgress == 87 and yProgress == 90) oColour <= 3'b110;
                    if(xProgress == 88 and yProgress == 90) oColour <= 3'b100;
                    if(xProgress == 89 and yProgress == 90) oColour <= 3'b111;
                    if(xProgress == 91 and yProgress == 90) oColour <= 3'b000;
                    if(xProgress == 69 and yProgress == 91) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 91) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 91) oColour <= 3'b110;
                    if(xProgress == 74 and yProgress == 91) oColour <= 3'b111;
                    if(xProgress == 75 and yProgress == 91) oColour <= 3'b110;
                    if(xProgress == 82 and yProgress == 91) oColour <= 3'b100;
                    if(xProgress == 83 and yProgress == 91) oColour <= 3'b110;
                    if(xProgress == 86 and yProgress == 91) oColour <= 3'b100;
                    if(xProgress == 87 and yProgress == 91) oColour <= 3'b110;
                    if(xProgress == 89 and yProgress == 91) oColour <= 3'b100;
                    if(xProgress == 90 and yProgress == 91) oColour <= 3'b111;
                    if(xProgress == 93 and yProgress == 91) oColour <= 3'b000;
                    if(xProgress == 12 and yProgress == 92) oColour <= 3'b001;
                    if(xProgress == 13 and yProgress == 92) oColour <= 3'b000;
                    if(xProgress == 68 and yProgress == 92) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 92) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 92) oColour <= 3'b110;
                    if(xProgress == 77 and yProgress == 92) oColour <= 3'b100;
                    if(xProgress == 80 and yProgress == 92) oColour <= 3'b110;
                    if(xProgress == 82 and yProgress == 92) oColour <= 3'b100;
                    if(xProgress == 83 and yProgress == 92) oColour <= 3'b110;
                    if(xProgress == 86 and yProgress == 92) oColour <= 3'b100;
                    if(xProgress == 88 and yProgress == 92) oColour <= 3'b110;
                    if(xProgress == 89 and yProgress == 92) oColour <= 3'b100;
                    if(xProgress == 90 and yProgress == 92) oColour <= 3'b111;
                    if(xProgress == 94 and yProgress == 92) oColour <= 3'b000;
                    if(xProgress == 67 and yProgress == 93) oColour <= 3'b111;
                    if(xProgress == 70 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 93) oColour <= 3'b110;
                    if(xProgress == 76 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 78 and yProgress == 93) oColour <= 3'b110;
                    if(xProgress == 79 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 80 and yProgress == 93) oColour <= 3'b110;
                    if(xProgress == 82 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 84 and yProgress == 93) oColour <= 3'b110;
                    if(xProgress == 87 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 88 and yProgress == 93) oColour <= 3'b110;
                    if(xProgress == 89 and yProgress == 93) oColour <= 3'b100;
                    if(xProgress == 92 and yProgress == 93) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 93) oColour <= 3'b000;
                    if(xProgress == 67 and yProgress == 94) oColour <= 3'b111;
                    if(xProgress == 69 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 70 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 71 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 72 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 73 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 75 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 76 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 77 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 79 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 80 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 83 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 84 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 87 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 88 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 89 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 90 and yProgress == 94) oColour <= 3'b110;
                    if(xProgress == 91 and yProgress == 94) oColour <= 3'b100;
                    if(xProgress == 93 and yProgress == 94) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 94) oColour <= 3'b000;
                    if(xProgress == 67 and yProgress == 95) oColour <= 3'b111;
                    if(xProgress == 69 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 70 and yProgress == 95) oColour <= 3'b110;
                    if(xProgress == 71 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 73 and yProgress == 95) oColour <= 3'b110;
                    if(xProgress == 75 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 80 and yProgress == 95) oColour <= 3'b110;
                    if(xProgress == 83 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 84 and yProgress == 95) oColour <= 3'b110;
                    if(xProgress == 87 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 89 and yProgress == 95) oColour <= 3'b110;
                    if(xProgress == 92 and yProgress == 95) oColour <= 3'b100;
                    if(xProgress == 93 and yProgress == 95) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 95) oColour <= 3'b000;
                    if(xProgress == 67 and yProgress == 96) oColour <= 3'b111;
                    if(xProgress == 70 and yProgress == 96) oColour <= 3'b100;
                    if(xProgress == 71 and yProgress == 96) oColour <= 3'b110;
                    if(xProgress == 73 and yProgress == 96) oColour <= 3'b100;
                    if(xProgress == 75 and yProgress == 96) oColour <= 3'b110;
                    if(xProgress == 77 and yProgress == 96) oColour <= 3'b100;
                    if(xProgress == 79 and yProgress == 96) oColour <= 3'b110;
                    if(xProgress == 80 and yProgress == 96) oColour <= 3'b100;
                    if(xProgress == 88 and yProgress == 96) oColour <= 3'b110;
                    if(xProgress == 92 and yProgress == 96) oColour <= 3'b100;
                    if(xProgress == 93 and yProgress == 96) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 96) oColour <= 3'b000;
                    if(xProgress == 68 and yProgress == 97) oColour <= 3'b111;
                    if(xProgress == 71 and yProgress == 97) oColour <= 3'b100;
                    if(xProgress == 75 and yProgress == 97) oColour <= 3'b110;
                    if(xProgress == 91 and yProgress == 97) oColour <= 3'b100;
                    if(xProgress == 93 and yProgress == 97) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 97) oColour <= 3'b000;
                    if(xProgress == 69 and yProgress == 98) oColour <= 3'b111;
                    if(xProgress == 74 and yProgress == 98) oColour <= 3'b100;
                    if(xProgress == 77 and yProgress == 98) oColour <= 3'b110;
                    if(xProgress == 90 and yProgress == 98) oColour <= 3'b100;
                    if(xProgress == 92 and yProgress == 98) oColour <= 3'b111;
                    if(xProgress == 95 and yProgress == 98) oColour <= 3'b000;
                    if(xProgress == 70 and yProgress == 99) oColour <= 3'b111;
                    if(xProgress == 76 and yProgress == 99) oColour <= 3'b100;
                    if(xProgress == 91 and yProgress == 99) oColour <= 3'b111;
                    if(xProgress == 94 and yProgress == 99) oColour <= 3'b000;
                    if(xProgress == 73 and yProgress == 100) oColour <= 3'b111;
                    if(xProgress == 93 and yProgress == 100) oColour <= 3'b000;
                    if(xProgress == 75 and yProgress == 101) oColour <= 3'b111;
                    if(xProgress == 92 and yProgress == 101) oColour <= 3'b000;
                    if(xProgress == 6 and yProgress == 102) oColour <= 3'b101;
                    if(xProgress == 12 and yProgress == 102) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 103) oColour <= 3'b101;
                    if(xProgress == 14 and yProgress == 103) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 104) oColour <= 3'b101;
                    if(xProgress == 6 and yProgress == 104) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 104) oColour <= 3'b101;
                    if(xProgress == 16 and yProgress == 104) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 105) oColour <= 3'b101;
                    if(xProgress == 4 and yProgress == 105) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 105) oColour <= 3'b101;
                    if(xProgress == 16 and yProgress == 105) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 106) oColour <= 3'b101;
                    if(xProgress == 4 and yProgress == 106) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 106) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 106) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 107) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 107) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 107) oColour <= 3'b101;
                    if(xProgress == 11 and yProgress == 107) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 107) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 107) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 108) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 108) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 108) oColour <= 3'b101;
                    if(xProgress == 11 and yProgress == 108) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 108) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 108) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 109) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 109) oColour <= 3'b100;
                    if(xProgress == 5 and yProgress == 109) oColour <= 3'b101;
                    if(xProgress == 7 and yProgress == 109) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 109) oColour <= 3'b101;
                    if(xProgress == 13 and yProgress == 109) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 109) oColour <= 3'b101;
                    if(xProgress == 20 and yProgress == 109) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 110) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 110) oColour <= 3'b100;
                    if(xProgress == 5 and yProgress == 110) oColour <= 3'b101;
                    if(xProgress == 7 and yProgress == 110) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 110) oColour <= 3'b101;
                    if(xProgress == 13 and yProgress == 110) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 110) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 110) oColour <= 3'b111;
                    if(xProgress == 19 and yProgress == 110) oColour <= 3'b101;
                    if(xProgress == 20 and yProgress == 110) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 111) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 111) oColour <= 3'b100;
                    if(xProgress == 5 and yProgress == 111) oColour <= 3'b101;
                    if(xProgress == 7 and yProgress == 111) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 111) oColour <= 3'b101;
                    if(xProgress == 13 and yProgress == 111) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 111) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 111) oColour <= 3'b111;
                    if(xProgress == 19 and yProgress == 111) oColour <= 3'b101;
                    if(xProgress == 20 and yProgress == 111) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 112) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 112) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 112) oColour <= 3'b101;
                    if(xProgress == 11 and yProgress == 112) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 112) oColour <= 3'b101;
                    if(xProgress == 20 and yProgress == 112) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 113) oColour <= 3'b101;
                    if(xProgress == 3 and yProgress == 113) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 113) oColour <= 3'b101;
                    if(xProgress == 11 and yProgress == 113) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 113) oColour <= 3'b101;
                    if(xProgress == 0 and yProgress == 114) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 114) oColour <= 3'b101;
                    if(xProgress == 4 and yProgress == 114) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 114) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 114) oColour <= 3'b110;
                    if(xProgress == 0 and yProgress == 115) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 6 and yProgress == 115) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 17 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 20 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 24 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 27 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 28 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 31 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 32 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 35 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 36 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 39 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 40 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 43 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 44 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 47 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 48 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 51 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 52 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 55 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 56 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 59 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 60 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 63 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 64 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 67 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 68 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 71 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 72 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 75 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 76 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 79 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 80 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 83 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 84 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 87 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 88 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 91 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 92 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 95 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 96 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 99 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 100 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 103 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 104 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 107 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 108 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 111 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 112 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 115 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 116 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 119 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 120 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 123 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 124 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 127 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 128 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 131 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 132 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 135 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 136 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 139 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 140 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 143 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 144 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 147 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 148 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 151 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 152 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 155 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 156 and yProgress == 115) oColour <= 3'b110;
                    if(xProgress == 159 and yProgress == 115) oColour <= 3'b101;
                    if(xProgress == 0 and yProgress == 116) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 116) oColour <= 3'b101;
                    if(xProgress == 0 and yProgress == 117) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 117) oColour <= 3'b101;
                    if(xProgress == 16 and yProgress == 117) oColour <= 3'b000;
                end else
                if(selector = 2'b01) begin
                    if(xProgress == 0 and yProgress == 0) oColour <= 3'b000;
                    if(xProgress == 11 and yProgress == 2) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 2) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 3) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 3) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 3) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 3) oColour <= 3'b000;
                    if(xProgress == 8 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 10 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 4) oColour <= 3'b000;
                    if(xProgress == 7 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 12 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 19 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 5) oColour <= 3'b000;
                    if(xProgress == 6 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 10 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 6) oColour <= 3'b111;
                    if(xProgress == 12 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 18 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 6) oColour <= 3'b000;
                    if(xProgress == 6 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 9 and yProgress == 7) oColour <= 3'b111;
                    if(xProgress == 11 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 7) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 8 and yProgress == 8) oColour <= 3'b111;
                    if(xProgress == 10 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 8) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 8 and yProgress == 9) oColour <= 3'b111;
                    if(xProgress == 9 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 9) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 10) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 11) oColour <= 3'b000;
                    if(xProgress == 3 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 4 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 5 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 7 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 12) oColour <= 3'b000;
                    if(xProgress == 3 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 4 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 5 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 9 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 13) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 5 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 7 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 13 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 14 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 14) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 15) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 15) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 15) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 15) oColour <= 3'b000;
                    if(xProgress == 8 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 16) oColour <= 3'b110;
                    if(xProgress == 24 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 16) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 25 and yProgress == 17) oColour <= 3'b000;
                end else
                if (selector == 2'b10) begin
                    if(xProgress == 0 and yProgress == 0) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 1) oColour <= 3'b110;
                    if(xProgress == 3 and yProgress == 1) oColour <= 3'b000;
                    if(xProgress == 27 and yProgress == 1) oColour <= 3'b110;
                    if(xProgress == 28 and yProgress == 1) oColour <= 3'b000;
                    if(xProgress == 3 and yProgress == 2) oColour <= 3'b110;
                    if(xProgress == 5 and yProgress == 2) oColour <= 3'b000;
                    if(xProgress == 11 and yProgress == 2) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 2) oColour <= 3'b000;
                    if(xProgress == 25 and yProgress == 2) oColour <= 3'b110;
                    if(xProgress == 27 and yProgress == 2) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 3) oColour <= 3'b110;
                    if(xProgress == 6 and yProgress == 3) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 3) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 3) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 3) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 3) oColour <= 3'b000;
                    if(xProgress == 24 and yProgress == 3) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 3) oColour <= 3'b000;
                    if(xProgress == 8 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 10 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 4) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 4) oColour <= 3'b000;
                    if(xProgress == 23 and yProgress == 4) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 4) oColour <= 3'b000;
                    if(xProgress == 7 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 12 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 19 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 5) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 5) oColour <= 3'b000;
                    if(xProgress == 29 and yProgress == 5) oColour <= 3'b110;
                    if(xProgress == 1 and yProgress == 6) oColour <= 3'b000;
                    if(xProgress == 6 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 10 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 6) oColour <= 3'b111;
                    if(xProgress == 12 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 15 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 18 and yProgress == 6) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 6) oColour <= 3'b000;
                    if(xProgress == 28 and yProgress == 6) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 6) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 3 and yProgress == 7) oColour <= 3'b000;
                    if(xProgress == 6 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 9 and yProgress == 7) oColour <= 3'b111;
                    if(xProgress == 11 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 16 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 20 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 7) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 7) oColour <= 3'b000;
                    if(xProgress == 26 and yProgress == 7) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 7) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 4 and yProgress == 8) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 8 and yProgress == 8) oColour <= 3'b111;
                    if(xProgress == 10 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 15 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 19 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 22 and yProgress == 8) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 8) oColour <= 3'b000;
                    if(xProgress == 26 and yProgress == 8) oColour <= 3'b110;
                    if(xProgress == 27 and yProgress == 8) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 8 and yProgress == 9) oColour <= 3'b111;
                    if(xProgress == 9 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 21 and yProgress == 9) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 9) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 9) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 17 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 20 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 10) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 10) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 10) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 3 and yProgress == 11) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 12 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 16 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 11) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 11) oColour <= 3'b000;
                    if(xProgress == 29 and yProgress == 11) oColour <= 3'b110;
                    if(xProgress == 2 and yProgress == 12) oColour <= 3'b000;
                    if(xProgress == 3 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 4 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 5 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 6 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 7 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 10 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 13 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 23 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 24 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 12) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 12) oColour <= 3'b000;
                    if(xProgress == 28 and yProgress == 12) oColour <= 3'b110;
                    if(xProgress == 1 and yProgress == 13) oColour <= 3'b000;
                    if(xProgress == 3 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 4 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 5 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 7 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 9 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 14 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 17 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 18 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 21 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 23 and yProgress == 13) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 13) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 13) oColour <= 3'b000;
                    if(xProgress == 4 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 5 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 7 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 11 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 13 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 14 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 22 and yProgress == 14) oColour <= 3'b110;
                    if(xProgress == 26 and yProgress == 14) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 14) oColour <= 3'b000;
                    if(xProgress == 5 and yProgress == 15) oColour <= 3'b100;
                    if(xProgress == 9 and yProgress == 15) oColour <= 3'b110;
                    if(xProgress == 25 and yProgress == 15) oColour <= 3'b100;
                    if(xProgress == 27 and yProgress == 15) oColour <= 3'b000;
                    if(xProgress == 2 and yProgress == 16) oColour <= 3'b110;
                    if(xProgress == 4 and yProgress == 16) oColour <= 3'b000;
                    if(xProgress == 8 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 11 and yProgress == 16) oColour <= 3'b110;
                    if(xProgress == 24 and yProgress == 16) oColour <= 3'b100;
                    if(xProgress == 26 and yProgress == 16) oColour <= 3'b000;
                    if(xProgress == 27 and yProgress == 16) oColour <= 3'b110;
                    if(xProgress == 29 and yProgress == 16) oColour <= 3'b000;
                    if(xProgress == 1 and yProgress == 17) oColour <= 3'b110;
                    if(xProgress == 3 and yProgress == 17) oColour <= 3'b000;
                    if(xProgress == 10 and yProgress == 17) oColour <= 3'b100;
                    if(xProgress == 25 and yProgress == 17) oColour <= 3'b000;
                    if(xProgress == 29 and yProgress == 17) oColour <= 3'b110;
                    if(xProgress == 1 and yProgress == 18) oColour <= 3'b000;
                end


            end else begin
                oDone <= 1; 
            end

    

        end else
        if (curState == ) begin//pick up here
            //before you say anything, I had a python script write this for me
            
        end else
        //if(selector)
    end
    




endmodule