module helper(iResetn,iPlotBox,iBlack,iColour,iLoadX,iXY_Coord,clk,oX,oY,oColour,oPlot,oDone);
    parameter X_SCREEN_PIXELS = 8'd160;
    parameter Y_SCREEN_PIXELS = 7'd120;
    input iResetn, iPlotBox, iBlack, iLoadX;
    input [2:0] iColour;
    input [6:0] iXY_Coord;
    input clk;
    output reg [7:0] oX;      //transformed coordinates 
    output reg [6:0] oY;
    output reg [2:0] oColour;     
    output reg oPlot;       
    output reg oDone;  


    localparam  RESET        = 3'd0,
                LOADING      = 3'd1,
                DRAW_GAME    = 3'd2,
                PLOT         = 3'd3
                G_STEADY     = 3'd4,
                G_HIT        = 3'd5,
                G_RESET      = 3'd6;
    
    reg [2:0] curState, nextState;
    reg [7:0] Xsize;            //upper bound of counter
    reg [6:0] Ysize;
    reg [7:0] xProgress;        //counter
    reg [6:0] yProgress;

    reg [2:0] oColour;

    reg [15:0] counter;

    reg [1:0] selector; //used to select colours
    

    /*
    (RESET) -> reset all variables
    (LOADING) -> Clears screen (minus tape measure)
                                                                                (out) (DRAW_GAME) -> draws full game screen
    (PLOT) -> Does the plotting
    (G_STEADY) -> waits for one of 3 buttons to go to next state
    (G_HIT) -> draws the hat that has been hit
    (G_RESET) -> Draws hat back to original

    iBlack = start

    iLoadX = hit1
    iPlotBox = hit2
    iResetn = resetn


    Selector:
    00 - draw base screen
    01 - draw hh no outline
    10 - draw hh 'hit'
    */

    colourSelect c0(.clk(clk), .xProgress(xProgress), .yProgress(yProgress), .selector(selector), .col(oColour)); //h&&les what colour should be outputted

    always@(*) begin
        case(curState)
        RESET: begin
            if(iBlack) nextState <= LOADING;
            //nextState <= iBlack ? LOADING ? RESET;
        end
        LOADING: 
            nextState <= oDone ? LOADING : PLOT;
        //DRAW_GAME:
            //nextState <= oDone ? G_STEADY : DRAW_GAME;
        //    nextState <= oDone ? LOADING: PLOT; //switches when nextState is released
        PLOT:
            if(selector == 2'b00) //after drawing main screen should go to steady
                nextState <= oDone ? G_STEADY : PLOT;
            else if(selector == 2'b01) //after drawing
                nextState <= oDone? G_RESET : PLOT;
            else if(selector <= 2'b10)
                nextState
        G_STEADY: begin
            if(iLoadX) nextState <= G_HIT;
            else if (iPlotBox) nextState <= G_HIT;
            else if(iResetn) nextState <= RESET;
        end
        G_HIT:   
            nextState = iPlotBox ? G_HIT : PLOT; //switches on negedge
        G_RESET: 
            nextState = oDone ? G_STEADY : G_RESET;
        endcase
    end

    always@(posedge clk) begin
        if(!iResetn) curState <= RESET;
        else curState <= nextState;

        if(curState == LOADING) begin //do something
            //drawing full screen so
            oDone <= 0;
            oPlot <= 1;  
            //oColour <= 3'b000; 
            Xsize <= X_SCREEN_PIXELS - 1;
            Ysize <= Y_SCREEN_PIXELS - 1;  
            oX <= 0;
            oY <= 0;
            xProgress <= 0;
            yProgress <= 0;
            selector <= 2'b00
        end 
        //else if (curState == DRAW_GAME) begin

        //end else
        else if(curState = PLOT) begin
            if (!oDone) begin
                oPlot <= 1;  
                //oColour <= oColour; 
                if (xProgress < Xsize) begin
                    oX <= oX + 1; 
                    xProgress <= xProgress + 1;  
                end else begin
                //if (xProgress == Xsize) begin
                    oX <= oX - xProgress;  
                    xProgress <= 0; 
                    if (yProgress < Ysize) begin
                        oY <= oY + 1;  
                        yProgress <= yProgress + 1; 
                    end
                end
                if (xProgress == Xsize && yProgress == Ysize) begin
                    oDone <= 1;  
                    oPlot <= 0;  
                    xSize <= 29; //xSize is for upper bound (these are now being set for hard-hat)
                    ySize <= 19;
                end
                //oColours from python script are assigned in other module
            end else begin
                oDone <= 1; 
            end
        end 
        else if (curState == G_STEADY) begin//pick up here
            if(iLoadX) begin//nextState <= G_HIT; (hit 1)
                //set vars for G_HIT
                selector <= 2'b10;
                oX <= 8'd47;
                oY <= 8'd15;
                oDone <= 1'b0;
                //oPlot <= 1'b1;
            end
            else if (iPlotBox) begin//nextState <= G_HIT; (hit 2)
                selector <= 2'b10;
                oX <= 8'd97;
                oY <= 7'd31;
                oDone <= 1'b0;
            end
            else if(iResetn) begin //nextState <= RESET;
                selector <= 2'b00;
                oX <=0;
                oY <= 0;
                oDone <=0;
            end
            
        end 
        else if(curState == G_HIT) begin
            //does anything need to be done here?

        end
        else if(curState == G_RESET) begin
            
        end
        //is there more that happens here?
    end
    




endmodule




module colourSelect(clk, xProgress, yProgress, selector, col)
    input clk;
    input reg [7:0] xProgress;
    input reg [6:0] yProgress;
    input reg [1:0] selector;

    output reg [2:0] col;
    always@(posedge clk) begin
        if(selector == 2'b00) begin //draw game screen
            if(xProgress == 0 && yProgress == 0) oColour <= 3'b000;
            else if(xProgress == 56 && yProgress == 13) oColour <= 3'b111;
            else if(xProgress == 63 && yProgress == 13) oColour <= 3'b000;
            else if(xProgress == 55 && yProgress == 14) oColour <= 3'b111;
            else if(xProgress == 67 && yProgress == 14) oColour <= 3'b000;
            else if(xProgress == 53 && yProgress == 15) oColour <= 3'b111;
            else if(xProgress == 57 && yProgress == 15) oColour <= 3'b100;
            else if(xProgress == 62 && yProgress == 15) oColour <= 3'b111;
            else if(xProgress == 68 && yProgress == 15) oColour <= 3'b000;
            else if(xProgress == 52 && yProgress == 16) oColour <= 3'b111;
            else if(xProgress == 56 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 58 && yProgress == 16) oColour <= 3'b110;
            else if(xProgress == 61 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 66 && yProgress == 16) oColour <= 3'b111;
            else if(xProgress == 69 && yProgress == 16) oColour <= 3'b000;
            else if(xProgress == 51 && yProgress == 17) oColour <= 3'b111;
            else if(xProgress == 54 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 56 && yProgress == 17) oColour <= 3'b110;
            else if(xProgress == 57 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 58 && yProgress == 17) oColour <= 3'b110;
            else if(xProgress == 62 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 63 && yProgress == 17) oColour <= 3'b110;
            else if(xProgress == 65 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 67 && yProgress == 17) oColour <= 3'b111;
            else if(xProgress == 69 && yProgress == 17) oColour <= 3'b000;
            else if(xProgress == 50 && yProgress == 18) oColour <= 3'b111;
            else if(xProgress == 53 && yProgress == 18) oColour <= 3'b100;
            else if(xProgress == 55 && yProgress == 18) oColour <= 3'b110;
            else if(xProgress == 56 && yProgress == 18) oColour <= 3'b100;
            else if(xProgress == 57 && yProgress == 18) oColour <= 3'b110;
            else if(xProgress == 58 && yProgress == 18) oColour <= 3'b100;
            else if(xProgress == 60 && yProgress == 18) oColour <= 3'b110;
            else if(xProgress == 63 && yProgress == 18) oColour <= 3'b100;
            else if(xProgress == 65 && yProgress == 18) oColour <= 3'b110;
            else if(xProgress == 66 && yProgress == 18) oColour <= 3'b100;
            else if(xProgress == 67 && yProgress == 18) oColour <= 3'b111;
            else if(xProgress == 70 && yProgress == 18) oColour <= 3'b000;
            else if(xProgress == 49 && yProgress == 19) oColour <= 3'b111;
            else if(xProgress == 52 && yProgress == 19) oColour <= 3'b100;
            else if(xProgress == 56 && yProgress == 19) oColour <= 3'b110;
            else if(xProgress == 57 && yProgress == 19) oColour <= 3'b111;
            else if(xProgress == 58 && yProgress == 19) oColour <= 3'b110;
            else if(xProgress == 59 && yProgress == 19) oColour <= 3'b100;
            else if(xProgress == 61 && yProgress == 19) oColour <= 3'b110;
            else if(xProgress == 64 && yProgress == 19) oColour <= 3'b100;
            else if(xProgress == 68 && yProgress == 19) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 19) oColour <= 3'b000;
            else if(xProgress == 49 && yProgress == 20) oColour <= 3'b111;
            else if(xProgress == 52 && yProgress == 20) oColour <= 3'b100;
            else if(xProgress == 53 && yProgress == 20) oColour <= 3'b110;
            else if(xProgress == 55 && yProgress == 20) oColour <= 3'b111;
            else if(xProgress == 57 && yProgress == 20) oColour <= 3'b110;
            else if(xProgress == 61 && yProgress == 20) oColour <= 3'b100;
            else if(xProgress == 62 && yProgress == 20) oColour <= 3'b110;
            else if(xProgress == 65 && yProgress == 20) oColour <= 3'b100;
            else if(xProgress == 66 && yProgress == 20) oColour <= 3'b110;
            else if(xProgress == 68 && yProgress == 20) oColour <= 3'b100;
            else if(xProgress == 69 && yProgress == 20) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 20) oColour <= 3'b000;
            else if(xProgress == 49 && yProgress == 21) oColour <= 3'b111;
            else if(xProgress == 51 && yProgress == 21) oColour <= 3'b100;
            else if(xProgress == 53 && yProgress == 21) oColour <= 3'b110;
            else if(xProgress == 54 && yProgress == 21) oColour <= 3'b111;
            else if(xProgress == 56 && yProgress == 21) oColour <= 3'b110;
            else if(xProgress == 61 && yProgress == 21) oColour <= 3'b100;
            else if(xProgress == 63 && yProgress == 21) oColour <= 3'b110;
            else if(xProgress == 65 && yProgress == 21) oColour <= 3'b100;
            else if(xProgress == 67 && yProgress == 21) oColour <= 3'b110;
            else if(xProgress == 68 && yProgress == 21) oColour <= 3'b100;
            else if(xProgress == 69 && yProgress == 21) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 21) oColour <= 3'b000;
            else if(xProgress == 49 && yProgress == 22) oColour <= 3'b111;
            else if(xProgress == 51 && yProgress == 22) oColour <= 3'b100;
            else if(xProgress == 52 && yProgress == 22) oColour <= 3'b110;
            else if(xProgress == 54 && yProgress == 22) oColour <= 3'b111;
            else if(xProgress == 55 && yProgress == 22) oColour <= 3'b110;
            else if(xProgress == 62 && yProgress == 22) oColour <= 3'b100;
            else if(xProgress == 63 && yProgress == 22) oColour <= 3'b110;
            else if(xProgress == 66 && yProgress == 22) oColour <= 3'b100;
            else if(xProgress == 67 && yProgress == 22) oColour <= 3'b110;
            else if(xProgress == 69 && yProgress == 22) oColour <= 3'b100;
            else if(xProgress == 70 && yProgress == 22) oColour <= 3'b111;
            else if(xProgress == 73 && yProgress == 22) oColour <= 3'b000;
            else if(xProgress == 48 && yProgress == 23) oColour <= 3'b111;
            else if(xProgress == 51 && yProgress == 23) oColour <= 3'b100;
            else if(xProgress == 52 && yProgress == 23) oColour <= 3'b110;
            else if(xProgress == 57 && yProgress == 23) oColour <= 3'b100;
            else if(xProgress == 60 && yProgress == 23) oColour <= 3'b110;
            else if(xProgress == 62 && yProgress == 23) oColour <= 3'b100;
            else if(xProgress == 63 && yProgress == 23) oColour <= 3'b110;
            else if(xProgress == 66 && yProgress == 23) oColour <= 3'b100;
            else if(xProgress == 68 && yProgress == 23) oColour <= 3'b110;
            else if(xProgress == 69 && yProgress == 23) oColour <= 3'b100;
            else if(xProgress == 70 && yProgress == 23) oColour <= 3'b111;
            else if(xProgress == 74 && yProgress == 23) oColour <= 3'b000;
            else if(xProgress == 47 && yProgress == 24) oColour <= 3'b111;
            else if(xProgress == 50 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 52 && yProgress == 24) oColour <= 3'b110;
            else if(xProgress == 56 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 58 && yProgress == 24) oColour <= 3'b110;
            else if(xProgress == 59 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 60 && yProgress == 24) oColour <= 3'b110;
            else if(xProgress == 62 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 64 && yProgress == 24) oColour <= 3'b110;
            else if(xProgress == 67 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 68 && yProgress == 24) oColour <= 3'b110;
            else if(xProgress == 69 && yProgress == 24) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 24) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 24) oColour <= 3'b000;
            else if(xProgress == 47 && yProgress == 25) oColour <= 3'b111;
            else if(xProgress == 49 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 50 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 51 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 52 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 53 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 55 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 56 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 57 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 59 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 60 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 63 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 64 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 67 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 68 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 69 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 70 && yProgress == 25) oColour <= 3'b110;
            else if(xProgress == 71 && yProgress == 25) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 25) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 25) oColour <= 3'b000;
            else if(xProgress == 47 && yProgress == 26) oColour <= 3'b111;
            else if(xProgress == 49 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 50 && yProgress == 26) oColour <= 3'b110;
            else if(xProgress == 51 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 53 && yProgress == 26) oColour <= 3'b110;
            else if(xProgress == 55 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 60 && yProgress == 26) oColour <= 3'b110;
            else if(xProgress == 63 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 64 && yProgress == 26) oColour <= 3'b110;
            else if(xProgress == 67 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 69 && yProgress == 26) oColour <= 3'b110;
            else if(xProgress == 72 && yProgress == 26) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 26) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 26) oColour <= 3'b000;
            else if(xProgress == 47 && yProgress == 27) oColour <= 3'b111;
            else if(xProgress == 50 && yProgress == 27) oColour <= 3'b100;
            else if(xProgress == 51 && yProgress == 27) oColour <= 3'b110;
            else if(xProgress == 53 && yProgress == 27) oColour <= 3'b100;
            else if(xProgress == 55 && yProgress == 27) oColour <= 3'b110;
            else if(xProgress == 57 && yProgress == 27) oColour <= 3'b100;
            else if(xProgress == 59 && yProgress == 27) oColour <= 3'b110;
            else if(xProgress == 60 && yProgress == 27) oColour <= 3'b100;
            else if(xProgress == 68 && yProgress == 27) oColour <= 3'b110;
            else if(xProgress == 72 && yProgress == 27) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 27) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 27) oColour <= 3'b000;
            else if(xProgress == 48 && yProgress == 28) oColour <= 3'b111;
            else if(xProgress == 51 && yProgress == 28) oColour <= 3'b100;
            else if(xProgress == 55 && yProgress == 28) oColour <= 3'b110;
            else if(xProgress == 71 && yProgress == 28) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 28) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 28) oColour <= 3'b000;
            else if(xProgress == 49 && yProgress == 29) oColour <= 3'b111;
            else if(xProgress == 54 && yProgress == 29) oColour <= 3'b100;
            else if(xProgress == 57 && yProgress == 29) oColour <= 3'b110;
            else if(xProgress == 70 && yProgress == 29) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 29) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 29) oColour <= 3'b000;
            else if(xProgress == 50 && yProgress == 30) oColour <= 3'b111;
            else if(xProgress == 56 && yProgress == 30) oColour <= 3'b100;
            else if(xProgress == 71 && yProgress == 30) oColour <= 3'b111;
            else if(xProgress == 74 && yProgress == 30) oColour <= 3'b000;
            else if(xProgress == 53 && yProgress == 31) oColour <= 3'b111;
            else if(xProgress == 73 && yProgress == 31) oColour <= 3'b000;
            else if(xProgress == 106 && yProgress == 31) oColour <= 3'b111;
            else if(xProgress == 113 && yProgress == 31) oColour <= 3'b000;
            else if(xProgress == 55 && yProgress == 32) oColour <= 3'b111;
            else if(xProgress == 72 && yProgress == 32) oColour <= 3'b000;
            else if(xProgress == 105 && yProgress == 32) oColour <= 3'b111;
            else if(xProgress == 117 && yProgress == 32) oColour <= 3'b000;
            else if(xProgress == 103 && yProgress == 33) oColour <= 3'b111;
            else if(xProgress == 107 && yProgress == 33) oColour <= 3'b100;
            else if(xProgress == 112 && yProgress == 33) oColour <= 3'b111;
            else if(xProgress == 118 && yProgress == 33) oColour <= 3'b000;
            else if(xProgress == 102 && yProgress == 34) oColour <= 3'b111;
            else if(xProgress == 106 && yProgress == 34) oColour <= 3'b100;
            else if(xProgress == 108 && yProgress == 34) oColour <= 3'b110;
            else if(xProgress == 111 && yProgress == 34) oColour <= 3'b100;
            else if(xProgress == 116 && yProgress == 34) oColour <= 3'b111;
            else if(xProgress == 119 && yProgress == 34) oColour <= 3'b000;
            else if(xProgress == 101 && yProgress == 35) oColour <= 3'b111;
            else if(xProgress == 104 && yProgress == 35) oColour <= 3'b100;
            else if(xProgress == 106 && yProgress == 35) oColour <= 3'b110;
            else if(xProgress == 107 && yProgress == 35) oColour <= 3'b100;
            else if(xProgress == 108 && yProgress == 35) oColour <= 3'b110;
            else if(xProgress == 112 && yProgress == 35) oColour <= 3'b100;
            else if(xProgress == 113 && yProgress == 35) oColour <= 3'b110;
            else if(xProgress == 115 && yProgress == 35) oColour <= 3'b100;
            else if(xProgress == 117 && yProgress == 35) oColour <= 3'b111;
            else if(xProgress == 119 && yProgress == 35) oColour <= 3'b000;
            else if(xProgress == 100 && yProgress == 36) oColour <= 3'b111;
            else if(xProgress == 103 && yProgress == 36) oColour <= 3'b100;
            else if(xProgress == 105 && yProgress == 36) oColour <= 3'b110;
            else if(xProgress == 106 && yProgress == 36) oColour <= 3'b100;
            else if(xProgress == 107 && yProgress == 36) oColour <= 3'b110;
            else if(xProgress == 108 && yProgress == 36) oColour <= 3'b100;
            else if(xProgress == 110 && yProgress == 36) oColour <= 3'b110;
            else if(xProgress == 113 && yProgress == 36) oColour <= 3'b100;
            else if(xProgress == 115 && yProgress == 36) oColour <= 3'b110;
            else if(xProgress == 116 && yProgress == 36) oColour <= 3'b100;
            else if(xProgress == 117 && yProgress == 36) oColour <= 3'b111;
            else if(xProgress == 120 && yProgress == 36) oColour <= 3'b000;
            else if(xProgress == 99 && yProgress == 37) oColour <= 3'b111;
            else if(xProgress == 102 && yProgress == 37) oColour <= 3'b100;
            else if(xProgress == 106 && yProgress == 37) oColour <= 3'b110;
            else if(xProgress == 107 && yProgress == 37) oColour <= 3'b111;
            else if(xProgress == 108 && yProgress == 37) oColour <= 3'b110;
            else if(xProgress == 109 && yProgress == 37) oColour <= 3'b100;
            else if(xProgress == 111 && yProgress == 37) oColour <= 3'b110;
            else if(xProgress == 114 && yProgress == 37) oColour <= 3'b100;
            else if(xProgress == 118 && yProgress == 37) oColour <= 3'b111;
            else if(xProgress == 121 && yProgress == 37) oColour <= 3'b000;
            else if(xProgress == 99 && yProgress == 38) oColour <= 3'b111;
            else if(xProgress == 102 && yProgress == 38) oColour <= 3'b100;
            else if(xProgress == 103 && yProgress == 38) oColour <= 3'b110;
            else if(xProgress == 105 && yProgress == 38) oColour <= 3'b111;
            else if(xProgress == 107 && yProgress == 38) oColour <= 3'b110;
            else if(xProgress == 111 && yProgress == 38) oColour <= 3'b100;
            else if(xProgress == 112 && yProgress == 38) oColour <= 3'b110;
            else if(xProgress == 115 && yProgress == 38) oColour <= 3'b100;
            else if(xProgress == 116 && yProgress == 38) oColour <= 3'b110;
            else if(xProgress == 118 && yProgress == 38) oColour <= 3'b100;
            else if(xProgress == 119 && yProgress == 38) oColour <= 3'b111;
            else if(xProgress == 121 && yProgress == 38) oColour <= 3'b000;
            else if(xProgress == 99 && yProgress == 39) oColour <= 3'b111;
            else if(xProgress == 101 && yProgress == 39) oColour <= 3'b100;
            else if(xProgress == 103 && yProgress == 39) oColour <= 3'b110;
            else if(xProgress == 104 && yProgress == 39) oColour <= 3'b111;
            else if(xProgress == 106 && yProgress == 39) oColour <= 3'b110;
            else if(xProgress == 111 && yProgress == 39) oColour <= 3'b100;
            else if(xProgress == 113 && yProgress == 39) oColour <= 3'b110;
            else if(xProgress == 115 && yProgress == 39) oColour <= 3'b100;
            else if(xProgress == 117 && yProgress == 39) oColour <= 3'b110;
            else if(xProgress == 118 && yProgress == 39) oColour <= 3'b100;
            else if(xProgress == 119 && yProgress == 39) oColour <= 3'b111;
            else if(xProgress == 121 && yProgress == 39) oColour <= 3'b000;
            else if(xProgress == 99 && yProgress == 40) oColour <= 3'b111;
            else if(xProgress == 101 && yProgress == 40) oColour <= 3'b100;
            else if(xProgress == 102 && yProgress == 40) oColour <= 3'b110;
            else if(xProgress == 104 && yProgress == 40) oColour <= 3'b111;
            else if(xProgress == 105 && yProgress == 40) oColour <= 3'b110;
            else if(xProgress == 112 && yProgress == 40) oColour <= 3'b100;
            else if(xProgress == 113 && yProgress == 40) oColour <= 3'b110;
            else if(xProgress == 116 && yProgress == 40) oColour <= 3'b100;
            else if(xProgress == 117 && yProgress == 40) oColour <= 3'b110;
            else if(xProgress == 119 && yProgress == 40) oColour <= 3'b100;
            else if(xProgress == 120 && yProgress == 40) oColour <= 3'b111;
            else if(xProgress == 123 && yProgress == 40) oColour <= 3'b000;
            else if(xProgress == 98 && yProgress == 41) oColour <= 3'b111;
            else if(xProgress == 101 && yProgress == 41) oColour <= 3'b100;
            else if(xProgress == 102 && yProgress == 41) oColour <= 3'b110;
            else if(xProgress == 107 && yProgress == 41) oColour <= 3'b100;
            else if(xProgress == 110 && yProgress == 41) oColour <= 3'b110;
            else if(xProgress == 112 && yProgress == 41) oColour <= 3'b100;
            else if(xProgress == 113 && yProgress == 41) oColour <= 3'b110;
            else if(xProgress == 116 && yProgress == 41) oColour <= 3'b100;
            else if(xProgress == 118 && yProgress == 41) oColour <= 3'b110;
            else if(xProgress == 119 && yProgress == 41) oColour <= 3'b100;
            else if(xProgress == 120 && yProgress == 41) oColour <= 3'b111;
            else if(xProgress == 124 && yProgress == 41) oColour <= 3'b000;
            else if(xProgress == 97 && yProgress == 42) oColour <= 3'b111;
            else if(xProgress == 100 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 102 && yProgress == 42) oColour <= 3'b110;
            else if(xProgress == 106 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 108 && yProgress == 42) oColour <= 3'b110;
            else if(xProgress == 109 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 110 && yProgress == 42) oColour <= 3'b110;
            else if(xProgress == 112 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 114 && yProgress == 42) oColour <= 3'b110;
            else if(xProgress == 117 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 118 && yProgress == 42) oColour <= 3'b110;
            else if(xProgress == 119 && yProgress == 42) oColour <= 3'b100;
            else if(xProgress == 122 && yProgress == 42) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 42) oColour <= 3'b000;
            else if(xProgress == 97 && yProgress == 43) oColour <= 3'b111;
            else if(xProgress == 99 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 100 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 101 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 102 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 103 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 105 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 106 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 107 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 109 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 110 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 113 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 114 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 117 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 118 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 119 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 120 && yProgress == 43) oColour <= 3'b110;
            else if(xProgress == 121 && yProgress == 43) oColour <= 3'b100;
            else if(xProgress == 123 && yProgress == 43) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 43) oColour <= 3'b000;
            else if(xProgress == 97 && yProgress == 44) oColour <= 3'b111;
            else if(xProgress == 99 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 100 && yProgress == 44) oColour <= 3'b110;
            else if(xProgress == 101 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 103 && yProgress == 44) oColour <= 3'b110;
            else if(xProgress == 105 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 110 && yProgress == 44) oColour <= 3'b110;
            else if(xProgress == 113 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 114 && yProgress == 44) oColour <= 3'b110;
            else if(xProgress == 117 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 119 && yProgress == 44) oColour <= 3'b110;
            else if(xProgress == 122 && yProgress == 44) oColour <= 3'b100;
            else if(xProgress == 123 && yProgress == 44) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 44) oColour <= 3'b000;
            else if(xProgress == 97 && yProgress == 45) oColour <= 3'b111;
            else if(xProgress == 100 && yProgress == 45) oColour <= 3'b100;
            else if(xProgress == 101 && yProgress == 45) oColour <= 3'b110;
            else if(xProgress == 103 && yProgress == 45) oColour <= 3'b100;
            else if(xProgress == 105 && yProgress == 45) oColour <= 3'b110;
            else if(xProgress == 107 && yProgress == 45) oColour <= 3'b100;
            else if(xProgress == 109 && yProgress == 45) oColour <= 3'b110;
            else if(xProgress == 110 && yProgress == 45) oColour <= 3'b100;
            else if(xProgress == 118 && yProgress == 45) oColour <= 3'b110;
            else if(xProgress == 122 && yProgress == 45) oColour <= 3'b100;
            else if(xProgress == 123 && yProgress == 45) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 45) oColour <= 3'b000;
            else if(xProgress == 98 && yProgress == 46) oColour <= 3'b111;
            else if(xProgress == 101 && yProgress == 46) oColour <= 3'b100;
            else if(xProgress == 105 && yProgress == 46) oColour <= 3'b110;
            else if(xProgress == 121 && yProgress == 46) oColour <= 3'b100;
            else if(xProgress == 123 && yProgress == 46) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 46) oColour <= 3'b000;
            else if(xProgress == 99 && yProgress == 47) oColour <= 3'b111;
            else if(xProgress == 104 && yProgress == 47) oColour <= 3'b100;
            else if(xProgress == 107 && yProgress == 47) oColour <= 3'b110;
            else if(xProgress == 120 && yProgress == 47) oColour <= 3'b100;
            else if(xProgress == 122 && yProgress == 47) oColour <= 3'b111;
            else if(xProgress == 125 && yProgress == 47) oColour <= 3'b000;
            else if(xProgress == 100 && yProgress == 48) oColour <= 3'b111;
            else if(xProgress == 106 && yProgress == 48) oColour <= 3'b100;
            else if(xProgress == 121 && yProgress == 48) oColour <= 3'b111;
            else if(xProgress == 124 && yProgress == 48) oColour <= 3'b000;
            else if(xProgress == 103 && yProgress == 49) oColour <= 3'b111;
            else if(xProgress == 123 && yProgress == 49) oColour <= 3'b000;
            else if(xProgress == 105 && yProgress == 50) oColour <= 3'b111;
            else if(xProgress == 122 && yProgress == 50) oColour <= 3'b000;
            else if(xProgress == 19 && yProgress == 53) oColour <= 3'b111;
            else if(xProgress == 26 && yProgress == 53) oColour <= 3'b000;
            else if(xProgress == 18 && yProgress == 54) oColour <= 3'b111;
            else if(xProgress == 30 && yProgress == 54) oColour <= 3'b000;
            else if(xProgress == 16 && yProgress == 55) oColour <= 3'b111;
            else if(xProgress == 20 && yProgress == 55) oColour <= 3'b100;
            else if(xProgress == 25 && yProgress == 55) oColour <= 3'b111;
            else if(xProgress == 31 && yProgress == 55) oColour <= 3'b000;
            else if(xProgress == 15 && yProgress == 56) oColour <= 3'b111;
            else if(xProgress == 19 && yProgress == 56) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 56) oColour <= 3'b110;
            else if(xProgress == 24 && yProgress == 56) oColour <= 3'b100;
            else if(xProgress == 29 && yProgress == 56) oColour <= 3'b111;
            else if(xProgress == 32 && yProgress == 56) oColour <= 3'b000;
            else if(xProgress == 14 && yProgress == 57) oColour <= 3'b111;
            else if(xProgress == 17 && yProgress == 57) oColour <= 3'b100;
            else if(xProgress == 19 && yProgress == 57) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 57) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 57) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 57) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 57) oColour <= 3'b110;
            else if(xProgress == 28 && yProgress == 57) oColour <= 3'b100;
            else if(xProgress == 30 && yProgress == 57) oColour <= 3'b111;
            else if(xProgress == 32 && yProgress == 57) oColour <= 3'b000;
            else if(xProgress == 13 && yProgress == 58) oColour <= 3'b111;
            else if(xProgress == 16 && yProgress == 58) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 58) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 58) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 58) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 58) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 58) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 58) oColour <= 3'b100;
            else if(xProgress == 28 && yProgress == 58) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 58) oColour <= 3'b100;
            else if(xProgress == 30 && yProgress == 58) oColour <= 3'b111;
            else if(xProgress == 33 && yProgress == 58) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 59) oColour <= 3'b111;
            else if(xProgress == 15 && yProgress == 59) oColour <= 3'b100;
            else if(xProgress == 19 && yProgress == 59) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 59) oColour <= 3'b111;
            else if(xProgress == 21 && yProgress == 59) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 59) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 59) oColour <= 3'b110;
            else if(xProgress == 27 && yProgress == 59) oColour <= 3'b100;
            else if(xProgress == 31 && yProgress == 59) oColour <= 3'b111;
            else if(xProgress == 34 && yProgress == 59) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 60) oColour <= 3'b111;
            else if(xProgress == 15 && yProgress == 60) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 60) oColour <= 3'b110;
            else if(xProgress == 18 && yProgress == 60) oColour <= 3'b111;
            else if(xProgress == 20 && yProgress == 60) oColour <= 3'b110;
            else if(xProgress == 24 && yProgress == 60) oColour <= 3'b100;
            else if(xProgress == 25 && yProgress == 60) oColour <= 3'b110;
            else if(xProgress == 28 && yProgress == 60) oColour <= 3'b100;
            else if(xProgress == 29 && yProgress == 60) oColour <= 3'b110;
            else if(xProgress == 31 && yProgress == 60) oColour <= 3'b100;
            else if(xProgress == 32 && yProgress == 60) oColour <= 3'b111;
            else if(xProgress == 34 && yProgress == 60) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 61) oColour <= 3'b111;
            else if(xProgress == 14 && yProgress == 61) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 61) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 61) oColour <= 3'b111;
            else if(xProgress == 19 && yProgress == 61) oColour <= 3'b110;
            else if(xProgress == 24 && yProgress == 61) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 61) oColour <= 3'b110;
            else if(xProgress == 28 && yProgress == 61) oColour <= 3'b100;
            else if(xProgress == 30 && yProgress == 61) oColour <= 3'b110;
            else if(xProgress == 31 && yProgress == 61) oColour <= 3'b100;
            else if(xProgress == 32 && yProgress == 61) oColour <= 3'b111;
            else if(xProgress == 34 && yProgress == 61) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 62) oColour <= 3'b111;
            else if(xProgress == 14 && yProgress == 62) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 62) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 62) oColour <= 3'b111;
            else if(xProgress == 18 && yProgress == 62) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 62) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 62) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 62) oColour <= 3'b100;
            else if(xProgress == 30 && yProgress == 62) oColour <= 3'b110;
            else if(xProgress == 32 && yProgress == 62) oColour <= 3'b100;
            else if(xProgress == 33 && yProgress == 62) oColour <= 3'b111;
            else if(xProgress == 36 && yProgress == 62) oColour <= 3'b000;
            else if(xProgress == 11 && yProgress == 63) oColour <= 3'b111;
            else if(xProgress == 14 && yProgress == 63) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 63) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 63) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 63) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 63) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 63) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 63) oColour <= 3'b100;
            else if(xProgress == 31 && yProgress == 63) oColour <= 3'b110;
            else if(xProgress == 32 && yProgress == 63) oColour <= 3'b100;
            else if(xProgress == 33 && yProgress == 63) oColour <= 3'b111;
            else if(xProgress == 37 && yProgress == 63) oColour <= 3'b000;
            else if(xProgress == 135 && yProgress == 63) oColour <= 3'b111;
            else if(xProgress == 142 && yProgress == 63) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 64) oColour <= 3'b111;
            else if(xProgress == 13 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 64) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 64) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 64) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 64) oColour <= 3'b110;
            else if(xProgress == 30 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 31 && yProgress == 64) oColour <= 3'b110;
            else if(xProgress == 32 && yProgress == 64) oColour <= 3'b100;
            else if(xProgress == 35 && yProgress == 64) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 64) oColour <= 3'b000;
            else if(xProgress == 134 && yProgress == 64) oColour <= 3'b111;
            else if(xProgress == 146 && yProgress == 64) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 65) oColour <= 3'b111;
            else if(xProgress == 12 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 13 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 14 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 30 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 31 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 32 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 33 && yProgress == 65) oColour <= 3'b110;
            else if(xProgress == 34 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 36 && yProgress == 65) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 65) oColour <= 3'b000;
            else if(xProgress == 132 && yProgress == 65) oColour <= 3'b111;
            else if(xProgress == 136 && yProgress == 65) oColour <= 3'b100;
            else if(xProgress == 141 && yProgress == 65) oColour <= 3'b111;
            else if(xProgress == 147 && yProgress == 65) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 66) oColour <= 3'b111;
            else if(xProgress == 12 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 13 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 14 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 18 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 30 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 32 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 35 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 36 && yProgress == 66) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 66) oColour <= 3'b000;
            else if(xProgress == 131 && yProgress == 66) oColour <= 3'b111;
            else if(xProgress == 135 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 137 && yProgress == 66) oColour <= 3'b110;
            else if(xProgress == 140 && yProgress == 66) oColour <= 3'b100;
            else if(xProgress == 145 && yProgress == 66) oColour <= 3'b111;
            else if(xProgress == 148 && yProgress == 66) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 67) oColour <= 3'b111;
            else if(xProgress == 13 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 31 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 35 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 36 && yProgress == 67) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 67) oColour <= 3'b000;
            else if(xProgress == 130 && yProgress == 67) oColour <= 3'b111;
            else if(xProgress == 133 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 135 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 136 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 137 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 141 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 142 && yProgress == 67) oColour <= 3'b110;
            else if(xProgress == 144 && yProgress == 67) oColour <= 3'b100;
            else if(xProgress == 146 && yProgress == 67) oColour <= 3'b111;
            else if(xProgress == 148 && yProgress == 67) oColour <= 3'b000;
            else if(xProgress == 11 && yProgress == 68) oColour <= 3'b111;
            else if(xProgress == 14 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 68) oColour <= 3'b110;
            else if(xProgress == 34 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 36 && yProgress == 68) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 68) oColour <= 3'b000;
            else if(xProgress == 129 && yProgress == 68) oColour <= 3'b111;
            else if(xProgress == 132 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 134 && yProgress == 68) oColour <= 3'b110;
            else if(xProgress == 135 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 136 && yProgress == 68) oColour <= 3'b110;
            else if(xProgress == 137 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 139 && yProgress == 68) oColour <= 3'b110;
            else if(xProgress == 142 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 144 && yProgress == 68) oColour <= 3'b110;
            else if(xProgress == 145 && yProgress == 68) oColour <= 3'b100;
            else if(xProgress == 146 && yProgress == 68) oColour <= 3'b111;
            else if(xProgress == 149 && yProgress == 68) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 69) oColour <= 3'b111;
            else if(xProgress == 17 && yProgress == 69) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 69) oColour <= 3'b110;
            else if(xProgress == 33 && yProgress == 69) oColour <= 3'b100;
            else if(xProgress == 35 && yProgress == 69) oColour <= 3'b111;
            else if(xProgress == 38 && yProgress == 69) oColour <= 3'b000;
            else if(xProgress == 128 && yProgress == 69) oColour <= 3'b111;
            else if(xProgress == 131 && yProgress == 69) oColour <= 3'b100;
            else if(xProgress == 135 && yProgress == 69) oColour <= 3'b110;
            else if(xProgress == 136 && yProgress == 69) oColour <= 3'b111;
            else if(xProgress == 137 && yProgress == 69) oColour <= 3'b110;
            else if(xProgress == 138 && yProgress == 69) oColour <= 3'b100;
            else if(xProgress == 140 && yProgress == 69) oColour <= 3'b110;
            else if(xProgress == 143 && yProgress == 69) oColour <= 3'b100;
            else if(xProgress == 147 && yProgress == 69) oColour <= 3'b111;
            else if(xProgress == 150 && yProgress == 69) oColour <= 3'b000;
            else if(xProgress == 13 && yProgress == 70) oColour <= 3'b111;
            else if(xProgress == 19 && yProgress == 70) oColour <= 3'b100;
            else if(xProgress == 34 && yProgress == 70) oColour <= 3'b111;
            else if(xProgress == 37 && yProgress == 70) oColour <= 3'b000;
            else if(xProgress == 128 && yProgress == 70) oColour <= 3'b111;
            else if(xProgress == 131 && yProgress == 70) oColour <= 3'b100;
            else if(xProgress == 132 && yProgress == 70) oColour <= 3'b110;
            else if(xProgress == 134 && yProgress == 70) oColour <= 3'b111;
            else if(xProgress == 136 && yProgress == 70) oColour <= 3'b110;
            else if(xProgress == 140 && yProgress == 70) oColour <= 3'b100;
            else if(xProgress == 141 && yProgress == 70) oColour <= 3'b110;
            else if(xProgress == 144 && yProgress == 70) oColour <= 3'b100;
            else if(xProgress == 145 && yProgress == 70) oColour <= 3'b110;
            else if(xProgress == 147 && yProgress == 70) oColour <= 3'b100;
            else if(xProgress == 148 && yProgress == 70) oColour <= 3'b111;
            else if(xProgress == 150 && yProgress == 70) oColour <= 3'b000;
            else if(xProgress == 16 && yProgress == 71) oColour <= 3'b111;
            else if(xProgress == 36 && yProgress == 71) oColour <= 3'b000;
            else if(xProgress == 128 && yProgress == 71) oColour <= 3'b111;
            else if(xProgress == 130 && yProgress == 71) oColour <= 3'b100;
            else if(xProgress == 132 && yProgress == 71) oColour <= 3'b110;
            else if(xProgress == 133 && yProgress == 71) oColour <= 3'b111;
            else if(xProgress == 135 && yProgress == 71) oColour <= 3'b110;
            else if(xProgress == 140 && yProgress == 71) oColour <= 3'b100;
            else if(xProgress == 142 && yProgress == 71) oColour <= 3'b110;
            else if(xProgress == 144 && yProgress == 71) oColour <= 3'b100;
            else if(xProgress == 146 && yProgress == 71) oColour <= 3'b110;
            else if(xProgress == 147 && yProgress == 71) oColour <= 3'b100;
            else if(xProgress == 148 && yProgress == 71) oColour <= 3'b111;
            else if(xProgress == 150 && yProgress == 71) oColour <= 3'b000;
            else if(xProgress == 18 && yProgress == 72) oColour <= 3'b111;
            else if(xProgress == 35 && yProgress == 72) oColour <= 3'b000;
            else if(xProgress == 128 && yProgress == 72) oColour <= 3'b111;
            else if(xProgress == 130 && yProgress == 72) oColour <= 3'b100;
            else if(xProgress == 131 && yProgress == 72) oColour <= 3'b110;
            else if(xProgress == 133 && yProgress == 72) oColour <= 3'b111;
            else if(xProgress == 134 && yProgress == 72) oColour <= 3'b110;
            else if(xProgress == 141 && yProgress == 72) oColour <= 3'b100;
            else if(xProgress == 142 && yProgress == 72) oColour <= 3'b110;
            else if(xProgress == 145 && yProgress == 72) oColour <= 3'b100;
            else if(xProgress == 146 && yProgress == 72) oColour <= 3'b110;
            else if(xProgress == 148 && yProgress == 72) oColour <= 3'b100;
            else if(xProgress == 149 && yProgress == 72) oColour <= 3'b111;
            else if(xProgress == 152 && yProgress == 72) oColour <= 3'b000;
            else if(xProgress == 127 && yProgress == 73) oColour <= 3'b111;
            else if(xProgress == 130 && yProgress == 73) oColour <= 3'b100;
            else if(xProgress == 131 && yProgress == 73) oColour <= 3'b110;
            else if(xProgress == 136 && yProgress == 73) oColour <= 3'b100;
            else if(xProgress == 139 && yProgress == 73) oColour <= 3'b110;
            else if(xProgress == 141 && yProgress == 73) oColour <= 3'b100;
            else if(xProgress == 142 && yProgress == 73) oColour <= 3'b110;
            else if(xProgress == 145 && yProgress == 73) oColour <= 3'b100;
            else if(xProgress == 147 && yProgress == 73) oColour <= 3'b110;
            else if(xProgress == 148 && yProgress == 73) oColour <= 3'b100;
            else if(xProgress == 149 && yProgress == 73) oColour <= 3'b111;
            else if(xProgress == 153 && yProgress == 73) oColour <= 3'b000;
            else if(xProgress == 126 && yProgress == 74) oColour <= 3'b111;
            else if(xProgress == 129 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 131 && yProgress == 74) oColour <= 3'b110;
            else if(xProgress == 135 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 137 && yProgress == 74) oColour <= 3'b110;
            else if(xProgress == 138 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 139 && yProgress == 74) oColour <= 3'b110;
            else if(xProgress == 141 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 143 && yProgress == 74) oColour <= 3'b110;
            else if(xProgress == 146 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 147 && yProgress == 74) oColour <= 3'b110;
            else if(xProgress == 148 && yProgress == 74) oColour <= 3'b100;
            else if(xProgress == 151 && yProgress == 74) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 74) oColour <= 3'b000;
            else if(xProgress == 126 && yProgress == 75) oColour <= 3'b111;
            else if(xProgress == 128 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 129 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 130 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 131 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 132 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 134 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 135 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 136 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 138 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 139 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 142 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 143 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 146 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 147 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 148 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 149 && yProgress == 75) oColour <= 3'b110;
            else if(xProgress == 150 && yProgress == 75) oColour <= 3'b100;
            else if(xProgress == 152 && yProgress == 75) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 75) oColour <= 3'b000;
            else if(xProgress == 126 && yProgress == 76) oColour <= 3'b111;
            else if(xProgress == 128 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 129 && yProgress == 76) oColour <= 3'b110;
            else if(xProgress == 130 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 132 && yProgress == 76) oColour <= 3'b110;
            else if(xProgress == 134 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 139 && yProgress == 76) oColour <= 3'b110;
            else if(xProgress == 142 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 143 && yProgress == 76) oColour <= 3'b110;
            else if(xProgress == 146 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 148 && yProgress == 76) oColour <= 3'b110;
            else if(xProgress == 151 && yProgress == 76) oColour <= 3'b100;
            else if(xProgress == 152 && yProgress == 76) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 76) oColour <= 3'b000;
            else if(xProgress == 126 && yProgress == 77) oColour <= 3'b111;
            else if(xProgress == 129 && yProgress == 77) oColour <= 3'b100;
            else if(xProgress == 130 && yProgress == 77) oColour <= 3'b110;
            else if(xProgress == 132 && yProgress == 77) oColour <= 3'b100;
            else if(xProgress == 134 && yProgress == 77) oColour <= 3'b110;
            else if(xProgress == 136 && yProgress == 77) oColour <= 3'b100;
            else if(xProgress == 138 && yProgress == 77) oColour <= 3'b110;
            else if(xProgress == 139 && yProgress == 77) oColour <= 3'b100;
            else if(xProgress == 147 && yProgress == 77) oColour <= 3'b110;
            else if(xProgress == 151 && yProgress == 77) oColour <= 3'b100;
            else if(xProgress == 152 && yProgress == 77) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 77) oColour <= 3'b000;
            else if(xProgress == 127 && yProgress == 78) oColour <= 3'b111;
            else if(xProgress == 130 && yProgress == 78) oColour <= 3'b100;
            else if(xProgress == 134 && yProgress == 78) oColour <= 3'b110;
            else if(xProgress == 150 && yProgress == 78) oColour <= 3'b100;
            else if(xProgress == 152 && yProgress == 78) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 78) oColour <= 3'b000;
            else if(xProgress == 128 && yProgress == 79) oColour <= 3'b111;
            else if(xProgress == 133 && yProgress == 79) oColour <= 3'b100;
            else if(xProgress == 136 && yProgress == 79) oColour <= 3'b110;
            else if(xProgress == 149 && yProgress == 79) oColour <= 3'b100;
            else if(xProgress == 151 && yProgress == 79) oColour <= 3'b111;
            else if(xProgress == 154 && yProgress == 79) oColour <= 3'b000;
            else if(xProgress == 129 && yProgress == 80) oColour <= 3'b111;
            else if(xProgress == 135 && yProgress == 80) oColour <= 3'b100;
            else if(xProgress == 150 && yProgress == 80) oColour <= 3'b111;
            else if(xProgress == 153 && yProgress == 80) oColour <= 3'b000;
            else if(xProgress == 132 && yProgress == 81) oColour <= 3'b111;
            else if(xProgress == 152 && yProgress == 81) oColour <= 3'b000;
            else if(xProgress == 76 && yProgress == 82) oColour <= 3'b111;
            else if(xProgress == 83 && yProgress == 82) oColour <= 3'b000;
            else if(xProgress == 134 && yProgress == 82) oColour <= 3'b111;
            else if(xProgress == 151 && yProgress == 82) oColour <= 3'b000;
            else if(xProgress == 75 && yProgress == 83) oColour <= 3'b111;
            else if(xProgress == 87 && yProgress == 83) oColour <= 3'b000;
            else if(xProgress == 73 && yProgress == 84) oColour <= 3'b111;
            else if(xProgress == 77 && yProgress == 84) oColour <= 3'b100;
            else if(xProgress == 82 && yProgress == 84) oColour <= 3'b111;
            else if(xProgress == 88 && yProgress == 84) oColour <= 3'b000;
            else if(xProgress == 72 && yProgress == 85) oColour <= 3'b111;
            else if(xProgress == 76 && yProgress == 85) oColour <= 3'b100;
            else if(xProgress == 78 && yProgress == 85) oColour <= 3'b110;
            else if(xProgress == 81 && yProgress == 85) oColour <= 3'b100;
            else if(xProgress == 86 && yProgress == 85) oColour <= 3'b111;
            else if(xProgress == 89 && yProgress == 85) oColour <= 3'b000;
            else if(xProgress == 71 && yProgress == 86) oColour <= 3'b111;
            else if(xProgress == 74 && yProgress == 86) oColour <= 3'b100;
            else if(xProgress == 76 && yProgress == 86) oColour <= 3'b110;
            else if(xProgress == 77 && yProgress == 86) oColour <= 3'b100;
            else if(xProgress == 78 && yProgress == 86) oColour <= 3'b110;
            else if(xProgress == 82 && yProgress == 86) oColour <= 3'b100;
            else if(xProgress == 83 && yProgress == 86) oColour <= 3'b110;
            else if(xProgress == 85 && yProgress == 86) oColour <= 3'b100;
            else if(xProgress == 87 && yProgress == 86) oColour <= 3'b111;
            else if(xProgress == 89 && yProgress == 86) oColour <= 3'b000;
            else if(xProgress == 70 && yProgress == 87) oColour <= 3'b111;
            else if(xProgress == 73 && yProgress == 87) oColour <= 3'b100;
            else if(xProgress == 75 && yProgress == 87) oColour <= 3'b110;
            else if(xProgress == 76 && yProgress == 87) oColour <= 3'b100;
            else if(xProgress == 77 && yProgress == 87) oColour <= 3'b110;
            else if(xProgress == 78 && yProgress == 87) oColour <= 3'b100;
            else if(xProgress == 80 && yProgress == 87) oColour <= 3'b110;
            else if(xProgress == 83 && yProgress == 87) oColour <= 3'b100;
            else if(xProgress == 85 && yProgress == 87) oColour <= 3'b110;
            else if(xProgress == 86 && yProgress == 87) oColour <= 3'b100;
            else if(xProgress == 87 && yProgress == 87) oColour <= 3'b111;
            else if(xProgress == 90 && yProgress == 87) oColour <= 3'b000;
            else if(xProgress == 69 && yProgress == 88) oColour <= 3'b111;
            else if(xProgress == 72 && yProgress == 88) oColour <= 3'b100;
            else if(xProgress == 76 && yProgress == 88) oColour <= 3'b110;
            else if(xProgress == 77 && yProgress == 88) oColour <= 3'b111;
            else if(xProgress == 78 && yProgress == 88) oColour <= 3'b110;
            else if(xProgress == 79 && yProgress == 88) oColour <= 3'b100;
            else if(xProgress == 81 && yProgress == 88) oColour <= 3'b110;
            else if(xProgress == 84 && yProgress == 88) oColour <= 3'b100;
            else if(xProgress == 88 && yProgress == 88) oColour <= 3'b111;
            else if(xProgress == 91 && yProgress == 88) oColour <= 3'b000;
            else if(xProgress == 69 && yProgress == 89) oColour <= 3'b111;
            else if(xProgress == 72 && yProgress == 89) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 89) oColour <= 3'b110;
            else if(xProgress == 75 && yProgress == 89) oColour <= 3'b111;
            else if(xProgress == 77 && yProgress == 89) oColour <= 3'b110;
            else if(xProgress == 81 && yProgress == 89) oColour <= 3'b100;
            else if(xProgress == 82 && yProgress == 89) oColour <= 3'b110;
            else if(xProgress == 85 && yProgress == 89) oColour <= 3'b100;
            else if(xProgress == 86 && yProgress == 89) oColour <= 3'b110;
            else if(xProgress == 88 && yProgress == 89) oColour <= 3'b100;
            else if(xProgress == 89 && yProgress == 89) oColour <= 3'b111;
            else if(xProgress == 91 && yProgress == 89) oColour <= 3'b000;
            else if(xProgress == 69 && yProgress == 90) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 90) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 90) oColour <= 3'b110;
            else if(xProgress == 74 && yProgress == 90) oColour <= 3'b111;
            else if(xProgress == 76 && yProgress == 90) oColour <= 3'b110;
            else if(xProgress == 81 && yProgress == 90) oColour <= 3'b100;
            else if(xProgress == 83 && yProgress == 90) oColour <= 3'b110;
            else if(xProgress == 85 && yProgress == 90) oColour <= 3'b100;
            else if(xProgress == 87 && yProgress == 90) oColour <= 3'b110;
            else if(xProgress == 88 && yProgress == 90) oColour <= 3'b100;
            else if(xProgress == 89 && yProgress == 90) oColour <= 3'b111;
            else if(xProgress == 91 && yProgress == 90) oColour <= 3'b000;
            else if(xProgress == 69 && yProgress == 91) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 91) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 91) oColour <= 3'b110;
            else if(xProgress == 74 && yProgress == 91) oColour <= 3'b111;
            else if(xProgress == 75 && yProgress == 91) oColour <= 3'b110;
            else if(xProgress == 82 && yProgress == 91) oColour <= 3'b100;
            else if(xProgress == 83 && yProgress == 91) oColour <= 3'b110;
            else if(xProgress == 86 && yProgress == 91) oColour <= 3'b100;
            else if(xProgress == 87 && yProgress == 91) oColour <= 3'b110;
            else if(xProgress == 89 && yProgress == 91) oColour <= 3'b100;
            else if(xProgress == 90 && yProgress == 91) oColour <= 3'b111;
            else if(xProgress == 93 && yProgress == 91) oColour <= 3'b000;
            else if(xProgress == 12 && yProgress == 92) oColour <= 3'b001;
            else if(xProgress == 13 && yProgress == 92) oColour <= 3'b000;
            else if(xProgress == 68 && yProgress == 92) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 92) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 92) oColour <= 3'b110;
            else if(xProgress == 77 && yProgress == 92) oColour <= 3'b100;
            else if(xProgress == 80 && yProgress == 92) oColour <= 3'b110;
            else if(xProgress == 82 && yProgress == 92) oColour <= 3'b100;
            else if(xProgress == 83 && yProgress == 92) oColour <= 3'b110;
            else if(xProgress == 86 && yProgress == 92) oColour <= 3'b100;
            else if(xProgress == 88 && yProgress == 92) oColour <= 3'b110;
            else if(xProgress == 89 && yProgress == 92) oColour <= 3'b100;
            else if(xProgress == 90 && yProgress == 92) oColour <= 3'b111;
            else if(xProgress == 94 && yProgress == 92) oColour <= 3'b000;
            else if(xProgress == 67 && yProgress == 93) oColour <= 3'b111;
            else if(xProgress == 70 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 93) oColour <= 3'b110;
            else if(xProgress == 76 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 78 && yProgress == 93) oColour <= 3'b110;
            else if(xProgress == 79 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 80 && yProgress == 93) oColour <= 3'b110;
            else if(xProgress == 82 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 84 && yProgress == 93) oColour <= 3'b110;
            else if(xProgress == 87 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 88 && yProgress == 93) oColour <= 3'b110;
            else if(xProgress == 89 && yProgress == 93) oColour <= 3'b100;
            else if(xProgress == 92 && yProgress == 93) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 93) oColour <= 3'b000;
            else if(xProgress == 67 && yProgress == 94) oColour <= 3'b111;
            else if(xProgress == 69 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 70 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 71 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 72 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 73 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 75 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 76 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 77 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 79 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 80 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 83 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 84 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 87 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 88 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 89 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 90 && yProgress == 94) oColour <= 3'b110;
            else if(xProgress == 91 && yProgress == 94) oColour <= 3'b100;
            else if(xProgress == 93 && yProgress == 94) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 94) oColour <= 3'b000;
            else if(xProgress == 67 && yProgress == 95) oColour <= 3'b111;
            else if(xProgress == 69 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 70 && yProgress == 95) oColour <= 3'b110;
            else if(xProgress == 71 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 73 && yProgress == 95) oColour <= 3'b110;
            else if(xProgress == 75 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 80 && yProgress == 95) oColour <= 3'b110;
            else if(xProgress == 83 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 84 && yProgress == 95) oColour <= 3'b110;
            else if(xProgress == 87 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 89 && yProgress == 95) oColour <= 3'b110;
            else if(xProgress == 92 && yProgress == 95) oColour <= 3'b100;
            else if(xProgress == 93 && yProgress == 95) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 95) oColour <= 3'b000;
            else if(xProgress == 67 && yProgress == 96) oColour <= 3'b111;
            else if(xProgress == 70 && yProgress == 96) oColour <= 3'b100;
            else if(xProgress == 71 && yProgress == 96) oColour <= 3'b110;
            else if(xProgress == 73 && yProgress == 96) oColour <= 3'b100;
            else if(xProgress == 75 && yProgress == 96) oColour <= 3'b110;
            else if(xProgress == 77 && yProgress == 96) oColour <= 3'b100;
            else if(xProgress == 79 && yProgress == 96) oColour <= 3'b110;
            else if(xProgress == 80 && yProgress == 96) oColour <= 3'b100;
            else if(xProgress == 88 && yProgress == 96) oColour <= 3'b110;
            else if(xProgress == 92 && yProgress == 96) oColour <= 3'b100;
            else if(xProgress == 93 && yProgress == 96) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 96) oColour <= 3'b000;
            else if(xProgress == 68 && yProgress == 97) oColour <= 3'b111;
            else if(xProgress == 71 && yProgress == 97) oColour <= 3'b100;
            else if(xProgress == 75 && yProgress == 97) oColour <= 3'b110;
            else if(xProgress == 91 && yProgress == 97) oColour <= 3'b100;
            else if(xProgress == 93 && yProgress == 97) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 97) oColour <= 3'b000;
            else if(xProgress == 69 && yProgress == 98) oColour <= 3'b111;
            else if(xProgress == 74 && yProgress == 98) oColour <= 3'b100;
            else if(xProgress == 77 && yProgress == 98) oColour <= 3'b110;
            else if(xProgress == 90 && yProgress == 98) oColour <= 3'b100;
            else if(xProgress == 92 && yProgress == 98) oColour <= 3'b111;
            else if(xProgress == 95 && yProgress == 98) oColour <= 3'b000;
            else if(xProgress == 70 && yProgress == 99) oColour <= 3'b111;
            else if(xProgress == 76 && yProgress == 99) oColour <= 3'b100;
            else if(xProgress == 91 && yProgress == 99) oColour <= 3'b111;
            else if(xProgress == 94 && yProgress == 99) oColour <= 3'b000;
            else if(xProgress == 73 && yProgress == 100) oColour <= 3'b111;
            else if(xProgress == 93 && yProgress == 100) oColour <= 3'b000;
            else if(xProgress == 75 && yProgress == 101) oColour <= 3'b111;
            else if(xProgress == 92 && yProgress == 101) oColour <= 3'b000;
            else if(xProgress == 6 && yProgress == 102) oColour <= 3'b101;
            else if(xProgress == 12 && yProgress == 102) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 103) oColour <= 3'b101;
            else if(xProgress == 14 && yProgress == 103) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 104) oColour <= 3'b101;
            else if(xProgress == 6 && yProgress == 104) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 104) oColour <= 3'b101;
            else if(xProgress == 16 && yProgress == 104) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 105) oColour <= 3'b101;
            else if(xProgress == 4 && yProgress == 105) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 105) oColour <= 3'b101;
            else if(xProgress == 16 && yProgress == 105) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 106) oColour <= 3'b101;
            else if(xProgress == 4 && yProgress == 106) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 106) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 106) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 107) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 107) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 107) oColour <= 3'b101;
            else if(xProgress == 11 && yProgress == 107) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 107) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 107) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 108) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 108) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 108) oColour <= 3'b101;
            else if(xProgress == 11 && yProgress == 108) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 108) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 108) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 109) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 109) oColour <= 3'b100;
            else if(xProgress == 5 && yProgress == 109) oColour <= 3'b101;
            else if(xProgress == 7 && yProgress == 109) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 109) oColour <= 3'b101;
            else if(xProgress == 13 && yProgress == 109) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 109) oColour <= 3'b101;
            else if(xProgress == 20 && yProgress == 109) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 110) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 110) oColour <= 3'b100;
            else if(xProgress == 5 && yProgress == 110) oColour <= 3'b101;
            else if(xProgress == 7 && yProgress == 110) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 110) oColour <= 3'b101;
            else if(xProgress == 13 && yProgress == 110) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 110) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 110) oColour <= 3'b111;
            else if(xProgress == 19 && yProgress == 110) oColour <= 3'b101;
            else if(xProgress == 20 && yProgress == 110) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 111) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 111) oColour <= 3'b100;
            else if(xProgress == 5 && yProgress == 111) oColour <= 3'b101;
            else if(xProgress == 7 && yProgress == 111) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 111) oColour <= 3'b101;
            else if(xProgress == 13 && yProgress == 111) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 111) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 111) oColour <= 3'b111;
            else if(xProgress == 19 && yProgress == 111) oColour <= 3'b101;
            else if(xProgress == 20 && yProgress == 111) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 112) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 112) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 112) oColour <= 3'b101;
            else if(xProgress == 11 && yProgress == 112) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 112) oColour <= 3'b101;
            else if(xProgress == 20 && yProgress == 112) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 113) oColour <= 3'b101;
            else if(xProgress == 3 && yProgress == 113) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 113) oColour <= 3'b101;
            else if(xProgress == 11 && yProgress == 113) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 113) oColour <= 3'b101;
            else if(xProgress == 0 && yProgress == 114) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 114) oColour <= 3'b101;
            else if(xProgress == 4 && yProgress == 114) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 114) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 114) oColour <= 3'b110;
            else if(xProgress == 0 && yProgress == 115) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 6 && yProgress == 115) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 17 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 20 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 24 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 27 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 28 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 31 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 32 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 35 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 36 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 39 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 40 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 43 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 44 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 47 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 48 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 51 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 52 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 55 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 56 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 59 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 60 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 63 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 64 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 67 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 68 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 71 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 72 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 75 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 76 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 79 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 80 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 83 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 84 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 87 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 88 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 91 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 92 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 95 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 96 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 99 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 100 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 103 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 104 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 107 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 108 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 111 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 112 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 115 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 116 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 119 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 120 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 123 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 124 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 127 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 128 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 131 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 132 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 135 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 136 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 139 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 140 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 143 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 144 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 147 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 148 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 151 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 152 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 155 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 156 && yProgress == 115) oColour <= 3'b110;
            else if(xProgress == 159 && yProgress == 115) oColour <= 3'b101;
            else if(xProgress == 0 && yProgress == 116) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 116) oColour <= 3'b101;
            else if(xProgress == 0 && yProgress == 117) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 117) oColour <= 3'b101;
            else if(xProgress == 16 && yProgress == 117) oColour <= 3'b000;
        end 
        else if(selector = 2'b01) begin //draw regular hat
            if(xProgress == 0 && yProgress == 0) oColour <= 3'b000;
            else if(xProgress == 11 && yProgress == 2) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 2) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 3) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 3) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 3) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 3) oColour <= 3'b000;
            else if(xProgress == 8 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 10 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 4) oColour <= 3'b000;
            else if(xProgress == 7 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 12 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 19 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 5) oColour <= 3'b000;
            else if(xProgress == 6 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 10 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 6) oColour <= 3'b111;
            else if(xProgress == 12 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 18 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 6) oColour <= 3'b000;
            else if(xProgress == 6 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 9 && yProgress == 7) oColour <= 3'b111;
            else if(xProgress == 11 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 7) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 8 && yProgress == 8) oColour <= 3'b111;
            else if(xProgress == 10 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 8) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 8 && yProgress == 9) oColour <= 3'b111;
            else if(xProgress == 9 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 9) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 10) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 11) oColour <= 3'b000;
            else if(xProgress == 3 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 4 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 5 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 7 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 12) oColour <= 3'b000;
            else if(xProgress == 3 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 4 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 5 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 9 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 13) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 5 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 7 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 13 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 14 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 14) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 15) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 15) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 15) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 15) oColour <= 3'b000;
            else if(xProgress == 8 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 16) oColour <= 3'b110;
            else if(xProgress == 24 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 16) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 25 && yProgress == 17) oColour <= 3'b000;
        end 
        else if (selector == 2'b10) begin  //colour selector for "hit" hat
            if(xProgress == 0 && yProgress == 0) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 1) oColour <= 3'b110;
            else if(xProgress == 3 && yProgress == 1) oColour <= 3'b000;
            else if(xProgress == 27 && yProgress == 1) oColour <= 3'b110;
            else if(xProgress == 28 && yProgress == 1) oColour <= 3'b000;
            else if(xProgress == 3 && yProgress == 2) oColour <= 3'b110;
            else if(xProgress == 5 && yProgress == 2) oColour <= 3'b000;
            else if(xProgress == 11 && yProgress == 2) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 2) oColour <= 3'b000;
            else if(xProgress == 25 && yProgress == 2) oColour <= 3'b110;
            else if(xProgress == 27 && yProgress == 2) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 3) oColour <= 3'b110;
            else if(xProgress == 6 && yProgress == 3) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 3) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 3) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 3) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 3) oColour <= 3'b000;
            else if(xProgress == 24 && yProgress == 3) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 3) oColour <= 3'b000;
            else if(xProgress == 8 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 10 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 4) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 4) oColour <= 3'b000;
            else if(xProgress == 23 && yProgress == 4) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 4) oColour <= 3'b000;
            else if(xProgress == 7 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 12 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 19 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 5) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 5) oColour <= 3'b000;
            else if(xProgress == 29 && yProgress == 5) oColour <= 3'b110;
            else if(xProgress == 1 && yProgress == 6) oColour <= 3'b000;
            else if(xProgress == 6 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 10 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 6) oColour <= 3'b111;
            else if(xProgress == 12 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 15 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 18 && yProgress == 6) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 6) oColour <= 3'b000;
            else if(xProgress == 28 && yProgress == 6) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 6) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 3 && yProgress == 7) oColour <= 3'b000;
            else if(xProgress == 6 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 9 && yProgress == 7) oColour <= 3'b111;
            else if(xProgress == 11 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 16 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 20 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 7) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 7) oColour <= 3'b000;
            else if(xProgress == 26 && yProgress == 7) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 7) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 4 && yProgress == 8) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 8 && yProgress == 8) oColour <= 3'b111;
            else if(xProgress == 10 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 15 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 19 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 22 && yProgress == 8) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 8) oColour <= 3'b000;
            else if(xProgress == 26 && yProgress == 8) oColour <= 3'b110;
            else if(xProgress == 27 && yProgress == 8) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 8 && yProgress == 9) oColour <= 3'b111;
            else if(xProgress == 9 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 21 && yProgress == 9) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 9) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 9) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 17 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 20 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 10) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 10) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 10) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 3 && yProgress == 11) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 12 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 16 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 11) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 11) oColour <= 3'b000;
            else if(xProgress == 29 && yProgress == 11) oColour <= 3'b110;
            else if(xProgress == 2 && yProgress == 12) oColour <= 3'b000;
            else if(xProgress == 3 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 4 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 5 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 6 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 7 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 10 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 13 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 23 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 24 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 12) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 12) oColour <= 3'b000;
            else if(xProgress == 28 && yProgress == 12) oColour <= 3'b110;
            else if(xProgress == 1 && yProgress == 13) oColour <= 3'b000;
            else if(xProgress == 3 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 4 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 5 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 7 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 9 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 14 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 17 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 18 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 21 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 23 && yProgress == 13) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 13) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 13) oColour <= 3'b000;
            else if(xProgress == 4 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 5 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 7 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 11 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 13 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 14 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 22 && yProgress == 14) oColour <= 3'b110;
            else if(xProgress == 26 && yProgress == 14) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 14) oColour <= 3'b000;
            else if(xProgress == 5 && yProgress == 15) oColour <= 3'b100;
            else if(xProgress == 9 && yProgress == 15) oColour <= 3'b110;
            else if(xProgress == 25 && yProgress == 15) oColour <= 3'b100;
            else if(xProgress == 27 && yProgress == 15) oColour <= 3'b000;
            else if(xProgress == 2 && yProgress == 16) oColour <= 3'b110;
            else if(xProgress == 4 && yProgress == 16) oColour <= 3'b000;
            else if(xProgress == 8 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 11 && yProgress == 16) oColour <= 3'b110;
            else if(xProgress == 24 && yProgress == 16) oColour <= 3'b100;
            else if(xProgress == 26 && yProgress == 16) oColour <= 3'b000;
            else if(xProgress == 27 && yProgress == 16) oColour <= 3'b110;
            else if(xProgress == 29 && yProgress == 16) oColour <= 3'b000;
            else if(xProgress == 1 && yProgress == 17) oColour <= 3'b110;
            else if(xProgress == 3 && yProgress == 17) oColour <= 3'b000;
            else if(xProgress == 10 && yProgress == 17) oColour <= 3'b100;
            else if(xProgress == 25 && yProgress == 17) oColour <= 3'b000;
            else if(xProgress == 29 && yProgress == 17) oColour <= 3'b110;
            else if(xProgress == 1 && yProgress == 18) oColour <= 3'b000;
        end
    end

endmodule

module part2(iResetn,iPlotBox,iBlack,iColour,iLoadX,iXY_Coord,iClock,oX,oY,oColour,oPlot,oDone);
   //specify input
   parameter X_SCREEN_PIXELS = 8'd160;
   parameter Y_SCREEN_PIXELS = 7'd120;
   input wire iResetn, iPlotBox, iBlack, iLoadX;
   input wire [2:0] iColour;
   input wire [6:0] iXY_Coord;
   input wire 	    iClock;
   output  [7:0] oX;       
   output  [6:0] oY;
   output  [2:0] oColour;     
   output  oPlot;       
   output  oDone;    

   helper u0(.iResetn(iResetn),.iPlotBox(iPlotBox),.iBlack(iBlack),
      .iColour(iColour), .iLoadX(iLoadX),.iXY_Coord(iXY_Coord),
      .clk(iClock),.oX(oX),.oY(oY), .oColour(oColour),
      .oPlot(oPlot),.oDone(oDone));
endmodule 