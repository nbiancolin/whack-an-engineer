module scoreKeeper (clock, scoreReset, moleHit, score);
    input clock;
    input scoreReset;
    input [2:0] hit;
    output reg [7:0] score;


endmodule